module tan_LUT(input [11:0] angle, output reg [23:0] ratio);

        always @(*) begin
                case(angle)
                        12'b000000000_000: ratio = 24'b00000000_0000000000000000;
                        12'b000000000_011: ratio = 24'b00000000_0000000110101100;
                        12'b000000000_110: ratio = 24'b00000000_0000001101011001;
                        12'b000000001_001: ratio = 24'b00000000_0000010100000110;
                        12'b000000001_100: ratio = 24'b00000000_0000011010110100;
                        12'b000000001_111: ratio = 24'b00000000_0000100001100001;
                        12'b000000010_010: ratio = 24'b00000000_0000101000001110;
                        12'b000000010_101: ratio = 24'b00000000_0000101110111100;
                        12'b000000011_000: ratio = 24'b00000000_0000110101101010;
                        12'b000000011_011: ratio = 24'b00000000_0000111100011000;
                        12'b000000011_110: ratio = 24'b00000000_0001000011000111;
                        12'b000000100_001: ratio = 24'b00000000_0001001001110110;
                        12'b000000100_100: ratio = 24'b00000000_0001010000100101;
                        12'b000000100_111: ratio = 24'b00000000_0001010111010101;
                        12'b000000101_010: ratio = 24'b00000000_0001011110000101;
                        12'b000000101_101: ratio = 24'b00000000_0001100100110110;
                        12'b000000110_000: ratio = 24'b00000000_0001101011101000;
                        12'b000000110_011: ratio = 24'b00000000_0001110010011010;
                        12'b000000110_110: ratio = 24'b00000000_0001111001001100;
                        12'b000000111_001: ratio = 24'b00000000_0001111111111111;
                        12'b000000111_100: ratio = 24'b00000000_0010000110110011;
                        12'b000000111_111: ratio = 24'b00000000_0010001101101000;
                        12'b000001000_010: ratio = 24'b00000000_0010010100011110;
                        12'b000001000_101: ratio = 24'b00000000_0010011011010100;
                        12'b000001001_000: ratio = 24'b00000000_0010100010001011;
                        12'b000001001_011: ratio = 24'b00000000_0010101001000100;
                        12'b000001001_110: ratio = 24'b00000000_0010101111111101;
                        12'b000001010_001: ratio = 24'b00000000_0010110110110111;
                        12'b000001010_100: ratio = 24'b00000000_0010111101110010;
                        12'b000001010_111: ratio = 24'b00000000_0011000100101110;
                        12'b000001011_010: ratio = 24'b00000000_0011001011101011;
                        12'b000001011_101: ratio = 24'b00000000_0011010010101010;
                        12'b000001100_000: ratio = 24'b00000000_0011011001101010;
                        12'b000001100_011: ratio = 24'b00000000_0011100000101011;
                        12'b000001100_110: ratio = 24'b00000000_0011100111101101;
                        12'b000001101_001: ratio = 24'b00000000_0011101110110000;
                        12'b000001101_100: ratio = 24'b00000000_0011110101110101;
                        12'b000001101_111: ratio = 24'b00000000_0011111100111100;
                        12'b000001110_010: ratio = 24'b00000000_0100000100000100;
                        12'b000001110_101: ratio = 24'b00000000_0100001011001101;
                        12'b000001111_000: ratio = 24'b00000000_0100010010011000;
                        12'b000001111_011: ratio = 24'b00000000_0100011001100100;
                        12'b000001111_110: ratio = 24'b00000000_0100100000110011;
                        12'b000010000_001: ratio = 24'b00000000_0100101000000010;
                        12'b000010000_100: ratio = 24'b00000000_0100101111010100;
                        12'b000010000_111: ratio = 24'b00000000_0100110110101000;
                        12'b000010001_010: ratio = 24'b00000000_0100111101111101;
                        12'b000010001_101: ratio = 24'b00000000_0101000101010100;
                        12'b000010010_000: ratio = 24'b00000000_0101001100101101;
                        12'b000010010_011: ratio = 24'b00000000_0101010100001001;
                        12'b000010010_110: ratio = 24'b00000000_0101011011100110;
                        12'b000010011_001: ratio = 24'b00000000_0101100011000101;
                        12'b000010011_100: ratio = 24'b00000000_0101101010100111;
                        12'b000010011_111: ratio = 24'b00000000_0101110010001011;
                        12'b000010100_010: ratio = 24'b00000000_0101111001110001;
                        12'b000010100_101: ratio = 24'b00000000_0110000001011010;
                        12'b000010101_000: ratio = 24'b00000000_0110001001000100;
                        12'b000010101_011: ratio = 24'b00000000_0110010000110010;
                        12'b000010101_110: ratio = 24'b00000000_0110011000100010;
                        12'b000010110_001: ratio = 24'b00000000_0110100000010100;
                        12'b000010110_100: ratio = 24'b00000000_0110101000001001;
                        12'b000010110_111: ratio = 24'b00000000_0110110000000001;
                        12'b000010111_010: ratio = 24'b00000000_0110110111111100;
                        12'b000010111_101: ratio = 24'b00000000_0110111111111010;
                        12'b000011000_000: ratio = 24'b00000000_0111000111111010;
                        12'b000011000_011: ratio = 24'b00000000_0111001111111101;
                        12'b000011000_110: ratio = 24'b00000000_0111011000000100;
                        12'b000011001_001: ratio = 24'b00000000_0111100000001110;
                        12'b000011001_100: ratio = 24'b00000000_0111101000011011;
                        12'b000011001_111: ratio = 24'b00000000_0111110000101011;
                        12'b000011010_010: ratio = 24'b00000000_0111111000111110;
                        12'b000011010_101: ratio = 24'b00000000_1000000001010101;
                        12'b000011011_000: ratio = 24'b00000000_1000001001110000;
                        12'b000011011_011: ratio = 24'b00000000_1000010010001110;
                        12'b000011011_110: ratio = 24'b00000000_1000011010110000;
                        12'b000011100_001: ratio = 24'b00000000_1000100011010101;
                        12'b000011100_100: ratio = 24'b00000000_1000101011111111;
                        12'b000011100_111: ratio = 24'b00000000_1000110100101100;
                        12'b000011101_010: ratio = 24'b00000000_1000111101011101;
                        12'b000011101_101: ratio = 24'b00000000_1001000110010011;
                        12'b000011110_000: ratio = 24'b00000000_1001001111001101;
                        12'b000011110_011: ratio = 24'b00000000_1001011000001011;
                        12'b000011110_110: ratio = 24'b00000000_1001100001001101;
                        12'b000011111_001: ratio = 24'b00000000_1001101010010100;
                        12'b000011111_100: ratio = 24'b00000000_1001110011100000;
                        12'b000011111_111: ratio = 24'b00000000_1001111100110000;
                        12'b000100000_010: ratio = 24'b00000000_1010000110000110;
                        12'b000100000_101: ratio = 24'b00000000_1010001111100000;
                        12'b000100001_000: ratio = 24'b00000000_1010011000111111;
                        12'b000100001_011: ratio = 24'b00000000_1010100010100100;
                        12'b000100001_110: ratio = 24'b00000000_1010101100001101;
                        12'b000100010_001: ratio = 24'b00000000_1010110101111100;
                        12'b000100010_100: ratio = 24'b00000000_1010111111110001;
                        12'b000100010_111: ratio = 24'b00000000_1011001001101100;
                        12'b000100011_010: ratio = 24'b00000000_1011010011101100;
                        12'b000100011_101: ratio = 24'b00000000_1011011101110010;
                        12'b000100100_000: ratio = 24'b00000000_1011100111111110;
                        12'b000100100_011: ratio = 24'b00000000_1011110010010001;
                        12'b000100100_110: ratio = 24'b00000000_1011111100101010;
                        12'b000100101_001: ratio = 24'b00000000_1100000111001001;
                        12'b000100101_100: ratio = 24'b00000000_1100010001101111;
                        12'b000100101_111: ratio = 24'b00000000_1100011100011100;
                        12'b000100110_010: ratio = 24'b00000000_1100100111010000;
                        12'b000100110_101: ratio = 24'b00000000_1100110010001011;
                        12'b000100111_000: ratio = 24'b00000000_1100111101001110;
                        12'b000100111_011: ratio = 24'b00000000_1101001000011000;
                        12'b000100111_110: ratio = 24'b00000000_1101010011101001;
                        12'b000101000_001: ratio = 24'b00000000_1101011111000011;
                        12'b000101000_100: ratio = 24'b00000000_1101101010100101;
                        12'b000101000_111: ratio = 24'b00000000_1101110110001111;
                        12'b000101001_010: ratio = 24'b00000000_1110000010000001;
                        12'b000101001_101: ratio = 24'b00000000_1110001101111100;
                        12'b000101010_000: ratio = 24'b00000000_1110011010000000;
                        12'b000101010_011: ratio = 24'b00000000_1110100110001110;
                        12'b000101010_110: ratio = 24'b00000000_1110110010100100;
                        12'b000101011_001: ratio = 24'b00000000_1110111111000101;
                        12'b000101011_100: ratio = 24'b00000000_1111001011101111;
                        12'b000101011_111: ratio = 24'b00000000_1111011000100011;
                        12'b000101100_010: ratio = 24'b00000000_1111100101100010;
                        12'b000101100_101: ratio = 24'b00000000_1111110010101011;
                        12'b000101101_000: ratio = 24'b00000001_0000000000000000;
                        12'b000101101_011: ratio = 24'b00000001_0000001101011111;
                        12'b000101101_110: ratio = 24'b00000001_0000011011001010;
                        12'b000101110_001: ratio = 24'b00000001_0000101001000001;
                        12'b000101110_100: ratio = 24'b00000001_0000110111000100;
                        12'b000101110_111: ratio = 24'b00000001_0001000101010100;
                        12'b000101111_010: ratio = 24'b00000001_0001010011110000;
                        12'b000101111_101: ratio = 24'b00000001_0001100010011001;
                        12'b000110000_000: ratio = 24'b00000001_0001110001010001;
                        12'b000110000_011: ratio = 24'b00000001_0010000000010110;
                        12'b000110000_110: ratio = 24'b00000001_0010001111101001;
                        12'b000110001_001: ratio = 24'b00000001_0010011111001011;
                        12'b000110001_100: ratio = 24'b00000001_0010101110111100;
                        12'b000110001_111: ratio = 24'b00000001_0010111110111101;
                        12'b000110010_010: ratio = 24'b00000001_0011001111001110;
                        12'b000110010_101: ratio = 24'b00000001_0011011111101111;
                        12'b000110011_000: ratio = 24'b00000001_0011110000100010;
                        12'b000110011_011: ratio = 24'b00000001_0100000001100110;
                        12'b000110011_110: ratio = 24'b00000001_0100010010111100;
                        12'b000110100_001: ratio = 24'b00000001_0100100100100100;
                        12'b000110100_100: ratio = 24'b00000001_0100110110100000;
                        12'b000110100_111: ratio = 24'b00000001_0101001000101111;
                        12'b000110101_010: ratio = 24'b00000001_0101011011010011;
                        12'b000110101_101: ratio = 24'b00000001_0101101110001100;
                        12'b000110110_000: ratio = 24'b00000001_0110000001011010;
                        12'b000110110_011: ratio = 24'b00000001_0110010100111111;
                        12'b000110110_110: ratio = 24'b00000001_0110101000111011;
                        12'b000110111_001: ratio = 24'b00000001_0110111101001111;
                        12'b000110111_100: ratio = 24'b00000001_0111010001111011;
                        12'b000110111_111: ratio = 24'b00000001_0111100111000001;
                        12'b000111000_010: ratio = 24'b00000001_0111111100100001;
                        12'b000111000_101: ratio = 24'b00000001_1000010010011100;
                        12'b000111001_000: ratio = 24'b00000001_1000101000110100;
                        12'b000111001_011: ratio = 24'b00000001_1000111111101001;
                        12'b000111001_110: ratio = 24'b00000001_1001010110111100;
                        12'b000111010_001: ratio = 24'b00000001_1001101110101110;
                        12'b000111010_100: ratio = 24'b00000001_1010000111000001;
                        12'b000111010_111: ratio = 24'b00000001_1010011111110101;
                        12'b000111011_010: ratio = 24'b00000001_1010111001001100;
                        12'b000111011_101: ratio = 24'b00000001_1011010011000111;
                        12'b000111100_000: ratio = 24'b00000001_1011101101100111;
                        12'b000111100_011: ratio = 24'b00000001_1100001000101111;
                        12'b000111100_110: ratio = 24'b00000001_1100100100011110;
                        12'b000111101_001: ratio = 24'b00000001_1101000000111000;
                        12'b000111101_100: ratio = 24'b00000001_1101011101111110;
                        12'b000111101_111: ratio = 24'b00000001_1101111011110001;
                        12'b000111110_010: ratio = 24'b00000001_1110011010010011;
                        12'b000111110_101: ratio = 24'b00000001_1110111001100110;
                        12'b000111111_000: ratio = 24'b00000001_1111011001101101;
                        12'b000111111_011: ratio = 24'b00000001_1111111010101001;
                        12'b000111111_110: ratio = 24'b00000010_0000011100011101;
                        12'b001000000_001: ratio = 24'b00000010_0000111111001100;
                        12'b001000000_100: ratio = 24'b00000010_0001100010110111;
                        12'b001000000_111: ratio = 24'b00000010_0010000111100001;
                        12'b001000001_010: ratio = 24'b00000010_0010101101001110;
                        12'b001000001_101: ratio = 24'b00000010_0011010100000001;
                        12'b001000010_000: ratio = 24'b00000010_0011111011111100;
                        12'b001000010_011: ratio = 24'b00000010_0100100101000011;
                        12'b001000010_110: ratio = 24'b00000010_0101001111011011;
                        12'b001000011_001: ratio = 24'b00000010_0101111011000110;
                        12'b001000011_100: ratio = 24'b00000010_0110101000001001;
                        12'b001000011_111: ratio = 24'b00000010_0111010110101001;
                        12'b001000100_010: ratio = 24'b00000010_1000000110101011;
                        12'b001000100_101: ratio = 24'b00000010_1000111000010011;
                        12'b001000101_000: ratio = 24'b00000010_1001101011100111;
                        12'b001000101_011: ratio = 24'b00000010_1010100000101100;
                        12'b001000101_110: ratio = 24'b00000010_1011010111101011;
                        12'b001000110_001: ratio = 24'b00000010_1100010000101000;
                        12'b001000110_100: ratio = 24'b00000010_1101001011101011;
                        12'b001000110_111: ratio = 24'b00000010_1110001000111101;
                        12'b001000111_010: ratio = 24'b00000010_1111001000100110;
                        12'b001000111_101: ratio = 24'b00000011_0000001010101111;
                        12'b001001000_000: ratio = 24'b00000011_0001001111100011;
                        12'b001001000_011: ratio = 24'b00000011_0010010111001011;
                        12'b001001000_110: ratio = 24'b00000011_0011100001110100;
                        12'b001001001_001: ratio = 24'b00000011_0100101111101011;
                        12'b001001001_100: ratio = 24'b00000011_0110000000111101;
                        12'b001001001_111: ratio = 24'b00000011_0111010101111011;
                        12'b001001010_010: ratio = 24'b00000011_1000101110110101;
                        12'b001001010_101: ratio = 24'b00000011_1010001011111101;
                        12'b001001011_000: ratio = 24'b00000011_1011101101100111;
                        12'b001001011_011: ratio = 24'b00000011_1101010100001011;
                        12'b001001011_110: ratio = 24'b00000011_1111000000000000;
                        12'b001001100_001: ratio = 24'b00000100_0000110001100011;
                        12'b001001100_100: ratio = 24'b00000100_0010101001010001;
                        12'b001001100_111: ratio = 24'b00000100_0100100111101100;
                        12'b001001101_010: ratio = 24'b00000100_0110101101011011;
                        12'b001001101_101: ratio = 24'b00000100_1000111011001000;
                        12'b001001110_000: ratio = 24'b00000100_1011010001100010;
                        12'b001001110_011: ratio = 24'b00000100_1101110001100000;
                        12'b001001110_110: ratio = 24'b00000101_0000011011111111;
                        12'b001001111_001: ratio = 24'b00000101_0011010010000101;
                        12'b001001111_100: ratio = 24'b00000101_0110010101000000;
                        12'b001001111_111: ratio = 24'b00000101_1001100110001101;
                        12'b001010000_010: ratio = 24'b00000101_1101000111010101;
                        12'b001010000_101: ratio = 24'b00000110_0000111010010001;
                        12'b001010001_000: ratio = 24'b00000110_0101000001010010;
                        12'b001010001_011: ratio = 24'b00000110_1001011110111101;
                        12'b001010001_110: ratio = 24'b00000110_1110010110011001;
                        12'b001010010_001: ratio = 24'b00000111_0011101011010010;
                        12'b001010010_100: ratio = 24'b00000111_1001100010000011;
                        12'b001010010_111: ratio = 24'b00001000_0000000000000001;
                        12'b001010011_010: ratio = 24'b00001000_0111001011101110;
                        12'b001010011_101: ratio = 24'b00001000_1111001101010000;
                        12'b001010100_000: ratio = 24'b00001001_1000001110101101;
                        12'b001010100_011: ratio = 24'b00001010_0010011100110110;
                        12'b001010100_110: ratio = 24'b00001010_1110001000000111;
                        12'b001010101_001: ratio = 24'b00001011_1011100101111111;
                        12'b001010101_100: ratio = 24'b00001100_1011010011001001;
                        12'b001010101_111: ratio = 24'b00001101_1101110110101010;
                        12'b001010110_010: ratio = 24'b00001111_0100000111001110;
                        12'b001010110_101: ratio = 24'b00010000_1111010011110110;
                        12'b001010111_000: ratio = 24'b00010011_0001010011000101;
                        12'b001010111_011: ratio = 24'b00010101_1100111111001010;
                        12'b001010111_110: ratio = 24'b00011001_0111001110100010;
                        12'b001011000_001: ratio = 24'b00011110_1000101111111101;
                        12'b001011000_100: ratio = 24'b00100110_0011000000111110;
                        12'b001011000_111: ratio = 24'b00110010_1110110001001100;
                        12'b001011001_010: ratio = 24'b01001100_0110001111010111;
                        12'b001011001_101: ratio = 24'b10011000_1100100101011100;
                        12'b001011010_000: ratio = -(24'b00000000_1111111111111111);
                        12'b001011010_011: ratio = -(24'b10011000_1100100101011011);
                        12'b001011010_110: ratio = -(24'b01001100_0110001111010111);
                        12'b001011011_001: ratio = -(24'b00110010_1110110001001100);
                        12'b001011011_100: ratio = -(24'b00100110_0011000000111110);
                        12'b001011011_111: ratio = -(24'b00011110_1000101111111101);
                        12'b001011100_010: ratio = -(24'b00011001_0111001110100010);
                        12'b001011100_101: ratio = -(24'b00010101_1100111111001010);
                        12'b001011101_000: ratio = -(24'b00010011_0001010011000101);
                        12'b001011101_011: ratio = -(24'b00010000_1111010011110110);
                        12'b001011101_110: ratio = -(24'b00001111_0100000111001110);
                        12'b001011110_001: ratio = -(24'b00001101_1101110110101010);
                        12'b001011110_100: ratio = -(24'b00001100_1011010011001001);
                        12'b001011110_111: ratio = -(24'b00001011_1011100101111111);
                        12'b001011111_010: ratio = -(24'b00001010_1110001000000111);
                        12'b001011111_101: ratio = -(24'b00001010_0010011100110110);
                        12'b001100000_000: ratio = -(24'b00001001_1000001110101101);
                        12'b001100000_011: ratio = -(24'b00001000_1111001101010000);
                        12'b001100000_110: ratio = -(24'b00001000_0111001011101110);
                        12'b001100001_001: ratio = -(24'b00001000_0000000000000001);
                        12'b001100001_100: ratio = -(24'b00000111_1001100010000011);
                        12'b001100001_111: ratio = -(24'b00000111_0011101011010010);
                        12'b001100010_010: ratio = -(24'b00000110_1110010110011001);
                        12'b001100010_101: ratio = -(24'b00000110_1001011110111101);
                        12'b001100011_000: ratio = -(24'b00000110_0101000001010010);
                        12'b001100011_011: ratio = -(24'b00000110_0000111010010001);
                        12'b001100011_110: ratio = -(24'b00000101_1101000111010101);
                        12'b001100100_001: ratio = -(24'b00000101_1001100110001101);
                        12'b001100100_100: ratio = -(24'b00000101_0110010101000000);
                        12'b001100100_111: ratio = -(24'b00000101_0011010010000101);
                        12'b001100101_010: ratio = -(24'b00000101_0000011011111111);
                        12'b001100101_101: ratio = -(24'b00000100_1101110001100000);
                        12'b001100110_000: ratio = -(24'b00000100_1011010001100010);
                        12'b001100110_011: ratio = -(24'b00000100_1000111011001000);
                        12'b001100110_110: ratio = -(24'b00000100_0110101101011011);
                        12'b001100111_001: ratio = -(24'b00000100_0100100111101100);
                        12'b001100111_100: ratio = -(24'b00000100_0010101001010001);
                        12'b001100111_111: ratio = -(24'b00000100_0000110001100011);
                        12'b001101000_010: ratio = -(24'b00000011_1111000000000000);
                        12'b001101000_101: ratio = -(24'b00000011_1101010100001011);
                        12'b001101001_000: ratio = -(24'b00000011_1011101101100111);
                        12'b001101001_011: ratio = -(24'b00000011_1010001011111101);
                        12'b001101001_110: ratio = -(24'b00000011_1000101110110101);
                        12'b001101010_001: ratio = -(24'b00000011_0111010101111011);
                        12'b001101010_100: ratio = -(24'b00000011_0110000000111101);
                        12'b001101010_111: ratio = -(24'b00000011_0100101111101011);
                        12'b001101011_010: ratio = -(24'b00000011_0011100001110100);
                        12'b001101011_101: ratio = -(24'b00000011_0010010111001011);
                        12'b001101100_000: ratio = -(24'b00000011_0001001111100011);
                        12'b001101100_011: ratio = -(24'b00000011_0000001010101111);
                        12'b001101100_110: ratio = -(24'b00000010_1111001000100110);
                        12'b001101101_001: ratio = -(24'b00000010_1110001000111101);
                        12'b001101101_100: ratio = -(24'b00000010_1101001011101011);
                        12'b001101101_111: ratio = -(24'b00000010_1100010000101000);
                        12'b001101110_010: ratio = -(24'b00000010_1011010111101011);
                        12'b001101110_101: ratio = -(24'b00000010_1010100000101100);
                        12'b001101111_000: ratio = -(24'b00000010_1001101011100111);
                        12'b001101111_011: ratio = -(24'b00000010_1000111000010011);
                        12'b001101111_110: ratio = -(24'b00000010_1000000110101011);
                        12'b001110000_001: ratio = -(24'b00000010_0111010110101001);
                        12'b001110000_100: ratio = -(24'b00000010_0110101000001001);
                        12'b001110000_111: ratio = -(24'b00000010_0101111011000110);
                        12'b001110001_010: ratio = -(24'b00000010_0101001111011011);
                        12'b001110001_101: ratio = -(24'b00000010_0100100101000011);
                        12'b001110010_000: ratio = -(24'b00000010_0011111011111100);
                        12'b001110010_011: ratio = -(24'b00000010_0011010100000001);
                        12'b001110010_110: ratio = -(24'b00000010_0010101101001110);
                        12'b001110011_001: ratio = -(24'b00000010_0010000111100001);
                        12'b001110011_100: ratio = -(24'b00000010_0001100010110111);
                        12'b001110011_111: ratio = -(24'b00000010_0000111111001100);
                        12'b001110100_010: ratio = -(24'b00000010_0000011100011101);
                        12'b001110100_101: ratio = -(24'b00000001_1111111010101001);
                        12'b001110101_000: ratio = -(24'b00000001_1111011001101101);
                        12'b001110101_011: ratio = -(24'b00000001_1110111001100110);
                        12'b001110101_110: ratio = -(24'b00000001_1110011010010011);
                        12'b001110110_001: ratio = -(24'b00000001_1101111011110001);
                        12'b001110110_100: ratio = -(24'b00000001_1101011101111110);
                        12'b001110110_111: ratio = -(24'b00000001_1101000000111000);
                        12'b001110111_010: ratio = -(24'b00000001_1100100100011110);
                        12'b001110111_101: ratio = -(24'b00000001_1100001000101111);
                        12'b001111000_000: ratio = -(24'b00000001_1011101101100111);
                        12'b001111000_011: ratio = -(24'b00000001_1011010011000111);
                        12'b001111000_110: ratio = -(24'b00000001_1010111001001100);
                        12'b001111001_001: ratio = -(24'b00000001_1010011111110101);
                        12'b001111001_100: ratio = -(24'b00000001_1010000111000001);
                        12'b001111001_111: ratio = -(24'b00000001_1001101110101110);
                        12'b001111010_010: ratio = -(24'b00000001_1001010110111100);
                        12'b001111010_101: ratio = -(24'b00000001_1000111111101001);
                        12'b001111011_000: ratio = -(24'b00000001_1000101000110100);
                        12'b001111011_011: ratio = -(24'b00000001_1000010010011100);
                        12'b001111011_110: ratio = -(24'b00000001_0111111100100001);
                        12'b001111100_001: ratio = -(24'b00000001_0111100111000001);
                        12'b001111100_100: ratio = -(24'b00000001_0111010001111011);
                        12'b001111100_111: ratio = -(24'b00000001_0110111101001111);
                        12'b001111101_010: ratio = -(24'b00000001_0110101000111011);
                        12'b001111101_101: ratio = -(24'b00000001_0110010100111111);
                        12'b001111110_000: ratio = -(24'b00000001_0110000001011010);
                        12'b001111110_011: ratio = -(24'b00000001_0101101110001100);
                        12'b001111110_110: ratio = -(24'b00000001_0101011011010011);
                        12'b001111111_001: ratio = -(24'b00000001_0101001000101111);
                        12'b001111111_100: ratio = -(24'b00000001_0100110110100000);
                        12'b001111111_111: ratio = -(24'b00000001_0100100100100100);
                        12'b010000000_010: ratio = -(24'b00000001_0100010010111100);
                        12'b010000000_101: ratio = -(24'b00000001_0100000001100110);
                        12'b010000001_000: ratio = -(24'b00000001_0011110000100010);
                        12'b010000001_011: ratio = -(24'b00000001_0011011111101111);
                        12'b010000001_110: ratio = -(24'b00000001_0011001111001110);
                        12'b010000010_001: ratio = -(24'b00000001_0010111110111101);
                        12'b010000010_100: ratio = -(24'b00000001_0010101110111100);
                        12'b010000010_111: ratio = -(24'b00000001_0010011111001011);
                        12'b010000011_010: ratio = -(24'b00000001_0010001111101001);
                        12'b010000011_101: ratio = -(24'b00000001_0010000000010110);
                        12'b010000100_000: ratio = -(24'b00000001_0001110001010001);
                        12'b010000100_011: ratio = -(24'b00000001_0001100010011001);
                        12'b010000100_110: ratio = -(24'b00000001_0001010011110000);
                        12'b010000101_001: ratio = -(24'b00000001_0001000101010100);
                        12'b010000101_100: ratio = -(24'b00000001_0000110111000100);
                        12'b010000101_111: ratio = -(24'b00000001_0000101001000001);
                        12'b010000110_010: ratio = -(24'b00000001_0000011011001010);
                        12'b010000110_101: ratio = -(24'b00000001_0000001101011111);
                        12'b010000111_000: ratio = -(24'b00000000_1111111111111111);
                        12'b010000111_011: ratio = -(24'b00000000_1111110010101011);
                        12'b010000111_110: ratio = -(24'b00000000_1111100101100010);
                        12'b010001000_001: ratio = -(24'b00000000_1111011000100011);
                        12'b010001000_100: ratio = -(24'b00000000_1111001011101111);
                        12'b010001000_111: ratio = -(24'b00000000_1110111111000101);
                        12'b010001001_010: ratio = -(24'b00000000_1110110010100100);
                        12'b010001001_101: ratio = -(24'b00000000_1110100110001110);
                        12'b010001010_000: ratio = -(24'b00000000_1110011010000000);
                        12'b010001010_011: ratio = -(24'b00000000_1110001101111100);
                        12'b010001010_110: ratio = -(24'b00000000_1110000010000001);
                        12'b010001011_001: ratio = -(24'b00000000_1101110110001111);
                        12'b010001011_100: ratio = -(24'b00000000_1101101010100101);
                        12'b010001011_111: ratio = -(24'b00000000_1101011111000011);
                        12'b010001100_010: ratio = -(24'b00000000_1101010011101001);
                        12'b010001100_101: ratio = -(24'b00000000_1101001000011000);
                        12'b010001101_000: ratio = -(24'b00000000_1100111101001110);
                        12'b010001101_011: ratio = -(24'b00000000_1100110010001011);
                        12'b010001101_110: ratio = -(24'b00000000_1100100111010000);
                        12'b010001110_001: ratio = -(24'b00000000_1100011100011100);
                        12'b010001110_100: ratio = -(24'b00000000_1100010001101111);
                        12'b010001110_111: ratio = -(24'b00000000_1100000111001001);
                        12'b010001111_010: ratio = -(24'b00000000_1011111100101010);
                        12'b010001111_101: ratio = -(24'b00000000_1011110010010001);
                        12'b010010000_000: ratio = -(24'b00000000_1011100111111110);
                        12'b010010000_011: ratio = -(24'b00000000_1011011101110010);
                        12'b010010000_110: ratio = -(24'b00000000_1011010011101100);
                        12'b010010001_001: ratio = -(24'b00000000_1011001001101100);
                        12'b010010001_100: ratio = -(24'b00000000_1010111111110001);
                        12'b010010001_111: ratio = -(24'b00000000_1010110101111100);
                        12'b010010010_010: ratio = -(24'b00000000_1010101100001101);
                        12'b010010010_101: ratio = -(24'b00000000_1010100010100100);
                        12'b010010011_000: ratio = -(24'b00000000_1010011000111111);
                        12'b010010011_011: ratio = -(24'b00000000_1010001111100000);
                        12'b010010011_110: ratio = -(24'b00000000_1010000110000110);
                        12'b010010100_001: ratio = -(24'b00000000_1001111100110000);
                        12'b010010100_100: ratio = -(24'b00000000_1001110011100000);
                        12'b010010100_111: ratio = -(24'b00000000_1001101010010100);
                        12'b010010101_010: ratio = -(24'b00000000_1001100001001101);
                        12'b010010101_101: ratio = -(24'b00000000_1001011000001011);
                        12'b010010110_000: ratio = -(24'b00000000_1001001111001101);
                        12'b010010110_011: ratio = -(24'b00000000_1001000110010011);
                        12'b010010110_110: ratio = -(24'b00000000_1000111101011101);
                        12'b010010111_001: ratio = -(24'b00000000_1000110100101100);
                        12'b010010111_100: ratio = -(24'b00000000_1000101011111111);
                        12'b010010111_111: ratio = -(24'b00000000_1000100011010101);
                        12'b010011000_010: ratio = -(24'b00000000_1000011010110000);
                        12'b010011000_101: ratio = -(24'b00000000_1000010010001110);
                        12'b010011001_000: ratio = -(24'b00000000_1000001001110000);
                        12'b010011001_011: ratio = -(24'b00000000_1000000001010101);
                        12'b010011001_110: ratio = -(24'b00000000_0111111000111110);
                        12'b010011010_001: ratio = -(24'b00000000_0111110000101011);
                        12'b010011010_100: ratio = -(24'b00000000_0111101000011011);
                        12'b010011010_111: ratio = -(24'b00000000_0111100000001110);
                        12'b010011011_010: ratio = -(24'b00000000_0111011000000100);
                        12'b010011011_101: ratio = -(24'b00000000_0111001111111101);
                        12'b010011100_000: ratio = -(24'b00000000_0111000111111010);
                        12'b010011100_011: ratio = -(24'b00000000_0110111111111010);
                        12'b010011100_110: ratio = -(24'b00000000_0110110111111100);
                        12'b010011101_001: ratio = -(24'b00000000_0110110000000001);
                        12'b010011101_100: ratio = -(24'b00000000_0110101000001001);
                        12'b010011101_111: ratio = -(24'b00000000_0110100000010100);
                        12'b010011110_010: ratio = -(24'b00000000_0110011000100010);
                        12'b010011110_101: ratio = -(24'b00000000_0110010000110010);
                        12'b010011111_000: ratio = -(24'b00000000_0110001001000100);
                        12'b010011111_011: ratio = -(24'b00000000_0110000001011010);
                        12'b010011111_110: ratio = -(24'b00000000_0101111001110001);
                        12'b010100000_001: ratio = -(24'b00000000_0101110010001011);
                        12'b010100000_100: ratio = -(24'b00000000_0101101010100111);
                        12'b010100000_111: ratio = -(24'b00000000_0101100011000101);
                        12'b010100001_010: ratio = -(24'b00000000_0101011011100110);
                        12'b010100001_101: ratio = -(24'b00000000_0101010100001001);
                        12'b010100010_000: ratio = -(24'b00000000_0101001100101101);
                        12'b010100010_011: ratio = -(24'b00000000_0101000101010100);
                        12'b010100010_110: ratio = -(24'b00000000_0100111101111101);
                        12'b010100011_001: ratio = -(24'b00000000_0100110110101000);
                        12'b010100011_100: ratio = -(24'b00000000_0100101111010100);
                        12'b010100011_111: ratio = -(24'b00000000_0100101000000010);
                        12'b010100100_010: ratio = -(24'b00000000_0100100000110011);
                        12'b010100100_101: ratio = -(24'b00000000_0100011001100100);
                        12'b010100101_000: ratio = -(24'b00000000_0100010010011000);
                        12'b010100101_011: ratio = -(24'b00000000_0100001011001101);
                        12'b010100101_110: ratio = -(24'b00000000_0100000100000100);
                        12'b010100110_001: ratio = -(24'b00000000_0011111100111100);
                        12'b010100110_100: ratio = -(24'b00000000_0011110101110101);
                        12'b010100110_111: ratio = -(24'b00000000_0011101110110000);
                        12'b010100111_010: ratio = -(24'b00000000_0011100111101101);
                        12'b010100111_101: ratio = -(24'b00000000_0011100000101011);
                        12'b010101000_000: ratio = -(24'b00000000_0011011001101010);
                        12'b010101000_011: ratio = -(24'b00000000_0011010010101010);
                        12'b010101000_110: ratio = -(24'b00000000_0011001011101011);
                        12'b010101001_001: ratio = -(24'b00000000_0011000100101110);
                        12'b010101001_100: ratio = -(24'b00000000_0010111101110010);
                        12'b010101001_111: ratio = -(24'b00000000_0010110110110111);
                        12'b010101010_010: ratio = -(24'b00000000_0010101111111101);
                        12'b010101010_101: ratio = -(24'b00000000_0010101001000100);
                        12'b010101011_000: ratio = -(24'b00000000_0010100010001011);
                        12'b010101011_011: ratio = -(24'b00000000_0010011011010100);
                        12'b010101011_110: ratio = -(24'b00000000_0010010100011110);
                        12'b010101100_001: ratio = -(24'b00000000_0010001101101000);
                        12'b010101100_100: ratio = -(24'b00000000_0010000110110011);
                        12'b010101100_111: ratio = -(24'b00000000_0001111111111111);
                        12'b010101101_010: ratio = -(24'b00000000_0001111001001100);
                        12'b010101101_101: ratio = -(24'b00000000_0001110010011010);
                        12'b010101110_000: ratio = -(24'b00000000_0001101011101000);
                        12'b010101110_011: ratio = -(24'b00000000_0001100100110110);
                        12'b010101110_110: ratio = -(24'b00000000_0001011110000101);
                        12'b010101111_001: ratio = -(24'b00000000_0001010111010101);
                        12'b010101111_100: ratio = -(24'b00000000_0001010000100101);
                        12'b010101111_111: ratio = -(24'b00000000_0001001001110110);
                        12'b010110000_010: ratio = -(24'b00000000_0001000011000111);
                        12'b010110000_101: ratio = -(24'b00000000_0000111100011000);
                        12'b010110001_000: ratio = -(24'b00000000_0000110101101010);
                        12'b010110001_011: ratio = -(24'b00000000_0000101110111100);
                        12'b010110001_110: ratio = -(24'b00000000_0000101000001110);
                        12'b010110010_001: ratio = -(24'b00000000_0000100001100001);
                        12'b010110010_100: ratio = -(24'b00000000_0000011010110100);
                        12'b010110010_111: ratio = -(24'b00000000_0000010100000110);
                        12'b010110011_010: ratio = -(24'b00000000_0000001101011001);
                        12'b010110011_101: ratio = -(24'b00000000_0000000110101100);
                        12'b010110100_000: ratio = 24'b00000000_0000000000000000;
                        12'b010110100_011: ratio = 24'b00000000_0000000110101100;
                        12'b010110100_110: ratio = 24'b00000000_0000001101011001;
                        12'b010110101_001: ratio = 24'b00000000_0000010100000110;
                        12'b010110101_100: ratio = 24'b00000000_0000011010110100;
                        12'b010110101_111: ratio = 24'b00000000_0000100001100001;
                        12'b010110110_010: ratio = 24'b00000000_0000101000001110;
                        12'b010110110_101: ratio = 24'b00000000_0000101110111100;
                        12'b010110111_000: ratio = 24'b00000000_0000110101101010;
                        12'b010110111_011: ratio = 24'b00000000_0000111100011000;
                        12'b010110111_110: ratio = 24'b00000000_0001000011000111;
                        12'b010111000_001: ratio = 24'b00000000_0001001001110110;
                        12'b010111000_100: ratio = 24'b00000000_0001010000100101;
                        12'b010111000_111: ratio = 24'b00000000_0001010111010101;
                        12'b010111001_010: ratio = 24'b00000000_0001011110000101;
                        12'b010111001_101: ratio = 24'b00000000_0001100100110110;
                        12'b010111010_000: ratio = 24'b00000000_0001101011101000;
                        12'b010111010_011: ratio = 24'b00000000_0001110010011010;
                        12'b010111010_110: ratio = 24'b00000000_0001111001001100;
                        12'b010111011_001: ratio = 24'b00000000_0001111111111111;
                        12'b010111011_100: ratio = 24'b00000000_0010000110110011;
                        12'b010111011_111: ratio = 24'b00000000_0010001101101000;
                        12'b010111100_010: ratio = 24'b00000000_0010010100011110;
                        12'b010111100_101: ratio = 24'b00000000_0010011011010100;
                        12'b010111101_000: ratio = 24'b00000000_0010100010001011;
                        12'b010111101_011: ratio = 24'b00000000_0010101001000100;
                        12'b010111101_110: ratio = 24'b00000000_0010101111111101;
                        12'b010111110_001: ratio = 24'b00000000_0010110110110111;
                        12'b010111110_100: ratio = 24'b00000000_0010111101110010;
                        12'b010111110_111: ratio = 24'b00000000_0011000100101110;
                        12'b010111111_010: ratio = 24'b00000000_0011001011101011;
                        12'b010111111_101: ratio = 24'b00000000_0011010010101010;
                        12'b011000000_000: ratio = 24'b00000000_0011011001101010;
                        12'b011000000_011: ratio = 24'b00000000_0011100000101011;
                        12'b011000000_110: ratio = 24'b00000000_0011100111101101;
                        12'b011000001_001: ratio = 24'b00000000_0011101110110000;
                        12'b011000001_100: ratio = 24'b00000000_0011110101110101;
                        12'b011000001_111: ratio = 24'b00000000_0011111100111100;
                        12'b011000010_010: ratio = 24'b00000000_0100000100000100;
                        12'b011000010_101: ratio = 24'b00000000_0100001011001101;
                        12'b011000011_000: ratio = 24'b00000000_0100010010011000;
                        12'b011000011_011: ratio = 24'b00000000_0100011001100100;
                        12'b011000011_110: ratio = 24'b00000000_0100100000110011;
                        12'b011000100_001: ratio = 24'b00000000_0100101000000010;
                        12'b011000100_100: ratio = 24'b00000000_0100101111010100;
                        12'b011000100_111: ratio = 24'b00000000_0100110110101000;
                        12'b011000101_010: ratio = 24'b00000000_0100111101111101;
                        12'b011000101_101: ratio = 24'b00000000_0101000101010100;
                        12'b011000110_000: ratio = 24'b00000000_0101001100101101;
                        12'b011000110_011: ratio = 24'b00000000_0101010100001001;
                        12'b011000110_110: ratio = 24'b00000000_0101011011100110;
                        12'b011000111_001: ratio = 24'b00000000_0101100011000101;
                        12'b011000111_100: ratio = 24'b00000000_0101101010100111;
                        12'b011000111_111: ratio = 24'b00000000_0101110010001011;
                        12'b011001000_010: ratio = 24'b00000000_0101111001110001;
                        12'b011001000_101: ratio = 24'b00000000_0110000001011010;
                        12'b011001001_000: ratio = 24'b00000000_0110001001000100;
                        12'b011001001_011: ratio = 24'b00000000_0110010000110010;
                        12'b011001001_110: ratio = 24'b00000000_0110011000100010;
                        12'b011001010_001: ratio = 24'b00000000_0110100000010100;
                        12'b011001010_100: ratio = 24'b00000000_0110101000001001;
                        12'b011001010_111: ratio = 24'b00000000_0110110000000001;
                        12'b011001011_010: ratio = 24'b00000000_0110110111111100;
                        12'b011001011_101: ratio = 24'b00000000_0110111111111010;
                        12'b011001100_000: ratio = 24'b00000000_0111000111111010;
                        12'b011001100_011: ratio = 24'b00000000_0111001111111101;
                        12'b011001100_110: ratio = 24'b00000000_0111011000000100;
                        12'b011001101_001: ratio = 24'b00000000_0111100000001110;
                        12'b011001101_100: ratio = 24'b00000000_0111101000011011;
                        12'b011001101_111: ratio = 24'b00000000_0111110000101011;
                        12'b011001110_010: ratio = 24'b00000000_0111111000111110;
                        12'b011001110_101: ratio = 24'b00000000_1000000001010101;
                        12'b011001111_000: ratio = 24'b00000000_1000001001110000;
                        12'b011001111_011: ratio = 24'b00000000_1000010010001110;
                        12'b011001111_110: ratio = 24'b00000000_1000011010110000;
                        12'b011010000_001: ratio = 24'b00000000_1000100011010101;
                        12'b011010000_100: ratio = 24'b00000000_1000101011111111;
                        12'b011010000_111: ratio = 24'b00000000_1000110100101100;
                        12'b011010001_010: ratio = 24'b00000000_1000111101011101;
                        12'b011010001_101: ratio = 24'b00000000_1001000110010011;
                        12'b011010010_000: ratio = 24'b00000000_1001001111001101;
                        12'b011010010_011: ratio = 24'b00000000_1001011000001011;
                        12'b011010010_110: ratio = 24'b00000000_1001100001001101;
                        12'b011010011_001: ratio = 24'b00000000_1001101010010100;
                        12'b011010011_100: ratio = 24'b00000000_1001110011100000;
                        12'b011010011_111: ratio = 24'b00000000_1001111100110000;
                        12'b011010100_010: ratio = 24'b00000000_1010000110000110;
                        12'b011010100_101: ratio = 24'b00000000_1010001111100000;
                        12'b011010101_000: ratio = 24'b00000000_1010011000111111;
                        12'b011010101_011: ratio = 24'b00000000_1010100010100100;
                        12'b011010101_110: ratio = 24'b00000000_1010101100001101;
                        12'b011010110_001: ratio = 24'b00000000_1010110101111100;
                        12'b011010110_100: ratio = 24'b00000000_1010111111110001;
                        12'b011010110_111: ratio = 24'b00000000_1011001001101100;
                        12'b011010111_010: ratio = 24'b00000000_1011010011101100;
                        12'b011010111_101: ratio = 24'b00000000_1011011101110010;
                        12'b011011000_000: ratio = 24'b00000000_1011100111111110;
                        12'b011011000_011: ratio = 24'b00000000_1011110010010001;
                        12'b011011000_110: ratio = 24'b00000000_1011111100101010;
                        12'b011011001_001: ratio = 24'b00000000_1100000111001001;
                        12'b011011001_100: ratio = 24'b00000000_1100010001101111;
                        12'b011011001_111: ratio = 24'b00000000_1100011100011100;
                        12'b011011010_010: ratio = 24'b00000000_1100100111010000;
                        12'b011011010_101: ratio = 24'b00000000_1100110010001011;
                        12'b011011011_000: ratio = 24'b00000000_1100111101001110;
                        12'b011011011_011: ratio = 24'b00000000_1101001000011000;
                        12'b011011011_110: ratio = 24'b00000000_1101010011101001;
                        12'b011011100_001: ratio = 24'b00000000_1101011111000011;
                        12'b011011100_100: ratio = 24'b00000000_1101101010100101;
                        12'b011011100_111: ratio = 24'b00000000_1101110110001111;
                        12'b011011101_010: ratio = 24'b00000000_1110000010000001;
                        12'b011011101_101: ratio = 24'b00000000_1110001101111100;
                        12'b011011110_000: ratio = 24'b00000000_1110011010000000;
                        12'b011011110_011: ratio = 24'b00000000_1110100110001110;
                        12'b011011110_110: ratio = 24'b00000000_1110110010100100;
                        12'b011011111_001: ratio = 24'b00000000_1110111111000101;
                        12'b011011111_100: ratio = 24'b00000000_1111001011101111;
                        12'b011011111_111: ratio = 24'b00000000_1111011000100011;
                        12'b011100000_010: ratio = 24'b00000000_1111100101100010;
                        12'b011100000_101: ratio = 24'b00000000_1111110010101011;
                        12'b011100001_000: ratio = 24'b00000001_0000000000000000;
                        12'b011100001_011: ratio = 24'b00000001_0000001101011111;
                        12'b011100001_110: ratio = 24'b00000001_0000011011001010;
                        12'b011100010_001: ratio = 24'b00000001_0000101001000001;
                        12'b011100010_100: ratio = 24'b00000001_0000110111000100;
                        12'b011100010_111: ratio = 24'b00000001_0001000101010100;
                        12'b011100011_010: ratio = 24'b00000001_0001010011110000;
                        12'b011100011_101: ratio = 24'b00000001_0001100010011001;
                        12'b011100100_000: ratio = 24'b00000001_0001110001010001;
                        12'b011100100_011: ratio = 24'b00000001_0010000000010110;
                        12'b011100100_110: ratio = 24'b00000001_0010001111101001;
                        12'b011100101_001: ratio = 24'b00000001_0010011111001011;
                        12'b011100101_100: ratio = 24'b00000001_0010101110111100;
                        12'b011100101_111: ratio = 24'b00000001_0010111110111101;
                        12'b011100110_010: ratio = 24'b00000001_0011001111001110;
                        12'b011100110_101: ratio = 24'b00000001_0011011111101111;
                        12'b011100111_000: ratio = 24'b00000001_0011110000100010;
                        12'b011100111_011: ratio = 24'b00000001_0100000001100110;
                        12'b011100111_110: ratio = 24'b00000001_0100010010111100;
                        12'b011101000_001: ratio = 24'b00000001_0100100100100100;
                        12'b011101000_100: ratio = 24'b00000001_0100110110100000;
                        12'b011101000_111: ratio = 24'b00000001_0101001000101111;
                        12'b011101001_010: ratio = 24'b00000001_0101011011010011;
                        12'b011101001_101: ratio = 24'b00000001_0101101110001100;
                        12'b011101010_000: ratio = 24'b00000001_0110000001011010;
                        12'b011101010_011: ratio = 24'b00000001_0110010100111111;
                        12'b011101010_110: ratio = 24'b00000001_0110101000111011;
                        12'b011101011_001: ratio = 24'b00000001_0110111101001111;
                        12'b011101011_100: ratio = 24'b00000001_0111010001111011;
                        12'b011101011_111: ratio = 24'b00000001_0111100111000001;
                        12'b011101100_010: ratio = 24'b00000001_0111111100100001;
                        12'b011101100_101: ratio = 24'b00000001_1000010010011100;
                        12'b011101101_000: ratio = 24'b00000001_1000101000110100;
                        12'b011101101_011: ratio = 24'b00000001_1000111111101001;
                        12'b011101101_110: ratio = 24'b00000001_1001010110111100;
                        12'b011101110_001: ratio = 24'b00000001_1001101110101110;
                        12'b011101110_100: ratio = 24'b00000001_1010000111000001;
                        12'b011101110_111: ratio = 24'b00000001_1010011111110101;
                        12'b011101111_010: ratio = 24'b00000001_1010111001001100;
                        12'b011101111_101: ratio = 24'b00000001_1011010011000111;
                        12'b011110000_000: ratio = 24'b00000001_1011101101100111;
                        12'b011110000_011: ratio = 24'b00000001_1100001000101111;
                        12'b011110000_110: ratio = 24'b00000001_1100100100011110;
                        12'b011110001_001: ratio = 24'b00000001_1101000000111000;
                        12'b011110001_100: ratio = 24'b00000001_1101011101111110;
                        12'b011110001_111: ratio = 24'b00000001_1101111011110001;
                        12'b011110010_010: ratio = 24'b00000001_1110011010010011;
                        12'b011110010_101: ratio = 24'b00000001_1110111001100110;
                        12'b011110011_000: ratio = 24'b00000001_1111011001101101;
                        12'b011110011_011: ratio = 24'b00000001_1111111010101001;
                        12'b011110011_110: ratio = 24'b00000010_0000011100011101;
                        12'b011110100_001: ratio = 24'b00000010_0000111111001100;
                        12'b011110100_100: ratio = 24'b00000010_0001100010110111;
                        12'b011110100_111: ratio = 24'b00000010_0010000111100001;
                        12'b011110101_010: ratio = 24'b00000010_0010101101001110;
                        12'b011110101_101: ratio = 24'b00000010_0011010100000001;
                        12'b011110110_000: ratio = 24'b00000010_0011111011111100;
                        12'b011110110_011: ratio = 24'b00000010_0100100101000011;
                        12'b011110110_110: ratio = 24'b00000010_0101001111011011;
                        12'b011110111_001: ratio = 24'b00000010_0101111011000110;
                        12'b011110111_100: ratio = 24'b00000010_0110101000001001;
                        12'b011110111_111: ratio = 24'b00000010_0111010110101001;
                        12'b011111000_010: ratio = 24'b00000010_1000000110101011;
                        12'b011111000_101: ratio = 24'b00000010_1000111000010011;
                        12'b011111001_000: ratio = 24'b00000010_1001101011100111;
                        12'b011111001_011: ratio = 24'b00000010_1010100000101100;
                        12'b011111001_110: ratio = 24'b00000010_1011010111101011;
                        12'b011111010_001: ratio = 24'b00000010_1100010000101000;
                        12'b011111010_100: ratio = 24'b00000010_1101001011101011;
                        12'b011111010_111: ratio = 24'b00000010_1110001000111101;
                        12'b011111011_010: ratio = 24'b00000010_1111001000100110;
                        12'b011111011_101: ratio = 24'b00000011_0000001010101111;
                        12'b011111100_000: ratio = 24'b00000011_0001001111100011;
                        12'b011111100_011: ratio = 24'b00000011_0010010111001011;
                        12'b011111100_110: ratio = 24'b00000011_0011100001110100;
                        12'b011111101_001: ratio = 24'b00000011_0100101111101011;
                        12'b011111101_100: ratio = 24'b00000011_0110000000111101;
                        12'b011111101_111: ratio = 24'b00000011_0111010101111011;
                        12'b011111110_010: ratio = 24'b00000011_1000101110110101;
                        12'b011111110_101: ratio = 24'b00000011_1010001011111101;
                        12'b011111111_000: ratio = 24'b00000011_1011101101100111;
                        12'b011111111_011: ratio = 24'b00000011_1101010100001011;
                        12'b011111111_110: ratio = 24'b00000011_1111000000000000;
                        12'b100000000_001: ratio = 24'b00000100_0000110001100011;
                        12'b100000000_100: ratio = 24'b00000100_0010101001010001;
                        12'b100000000_111: ratio = 24'b00000100_0100100111101100;
                        12'b100000001_010: ratio = 24'b00000100_0110101101011011;
                        12'b100000001_101: ratio = 24'b00000100_1000111011001000;
                        12'b100000010_000: ratio = 24'b00000100_1011010001100010;
                        12'b100000010_011: ratio = 24'b00000100_1101110001100000;
                        12'b100000010_110: ratio = 24'b00000101_0000011011111111;
                        12'b100000011_001: ratio = 24'b00000101_0011010010000101;
                        12'b100000011_100: ratio = 24'b00000101_0110010101000000;
                        12'b100000011_111: ratio = 24'b00000101_1001100110001101;
                        12'b100000100_010: ratio = 24'b00000101_1101000111010101;
                        12'b100000100_101: ratio = 24'b00000110_0000111010010001;
                        12'b100000101_000: ratio = 24'b00000110_0101000001010010;
                        12'b100000101_011: ratio = 24'b00000110_1001011110111101;
                        12'b100000101_110: ratio = 24'b00000110_1110010110011001;
                        12'b100000110_001: ratio = 24'b00000111_0011101011010010;
                        12'b100000110_100: ratio = 24'b00000111_1001100010000011;
                        12'b100000110_111: ratio = 24'b00001000_0000000000000001;
                        12'b100000111_010: ratio = 24'b00001000_0111001011101110;
                        12'b100000111_101: ratio = 24'b00001000_1111001101010000;
                        12'b100001000_000: ratio = 24'b00001001_1000001110101101;
                        12'b100001000_011: ratio = 24'b00001010_0010011100110110;
                        12'b100001000_110: ratio = 24'b00001010_1110001000000111;
                        12'b100001001_001: ratio = 24'b00001011_1011100101111111;
                        12'b100001001_100: ratio = 24'b00001100_1011010011001001;
                        12'b100001001_111: ratio = 24'b00001101_1101110110101010;
                        12'b100001010_010: ratio = 24'b00001111_0100000111001110;
                        12'b100001010_101: ratio = 24'b00010000_1111010011110110;
                        12'b100001011_000: ratio = 24'b00010011_0001010011000101;
                        12'b100001011_011: ratio = 24'b00010101_1100111111001010;
                        12'b100001011_110: ratio = 24'b00011001_0111001110100010;
                        12'b100001100_001: ratio = 24'b00011110_1000101111111101;
                        12'b100001100_100: ratio = 24'b00100110_0011000000111110;
                        12'b100001100_111: ratio = 24'b00110010_1110110001001100;
                        12'b100001101_010: ratio = 24'b01001100_0110001111010111;
                        12'b100001101_101: ratio = 24'b10011000_1100100101011101;
                        12'b100001110_000: ratio = -(24'b11111111_0000000000000000);
                        12'b100001110_011: ratio = -(24'b10011000_1100100101011011);
                        12'b100001110_110: ratio = -(24'b01001100_0110001111010111);
                        12'b100001111_001: ratio = -(24'b00110010_1110110001001100);
                        12'b100001111_100: ratio = -(24'b00100110_0011000000111110);
                        12'b100001111_111: ratio = -(24'b00011110_1000101111111101);
                        12'b100010000_010: ratio = -(24'b00011001_0111001110100010);
                        12'b100010000_101: ratio = -(24'b00010101_1100111111001010);
                        12'b100010001_000: ratio = -(24'b00010011_0001010011000101);
                        12'b100010001_011: ratio = -(24'b00010000_1111010011110110);
                        12'b100010001_110: ratio = -(24'b00001111_0100000111001110);
                        12'b100010010_001: ratio = -(24'b00001101_1101110110101010);
                        12'b100010010_100: ratio = -(24'b00001100_1011010011001001);
                        12'b100010010_111: ratio = -(24'b00001011_1011100101111111);
                        12'b100010011_010: ratio = -(24'b00001010_1110001000000111);
                        12'b100010011_101: ratio = -(24'b00001010_0010011100110110);
                        12'b100010100_000: ratio = -(24'b00001001_1000001110101101);
                        12'b100010100_011: ratio = -(24'b00001000_1111001101010000);
                        12'b100010100_110: ratio = -(24'b00001000_0111001011101110);
                        12'b100010101_001: ratio = -(24'b00001000_0000000000000001);
                        12'b100010101_100: ratio = -(24'b00000111_1001100010000011);
                        12'b100010101_111: ratio = -(24'b00000111_0011101011010010);
                        12'b100010110_010: ratio = -(24'b00000110_1110010110011001);
                        12'b100010110_101: ratio = -(24'b00000110_1001011110111101);
                        12'b100010111_000: ratio = -(24'b00000110_0101000001010010);
                        12'b100010111_011: ratio = -(24'b00000110_0000111010010001);
                        12'b100010111_110: ratio = -(24'b00000101_1101000111010101);
                        12'b100011000_001: ratio = -(24'b00000101_1001100110001101);
                        12'b100011000_100: ratio = -(24'b00000101_0110010101000000);
                        12'b100011000_111: ratio = -(24'b00000101_0011010010000101);
                        12'b100011001_010: ratio = -(24'b00000101_0000011011111111);
                        12'b100011001_101: ratio = -(24'b00000100_1101110001100000);
                        12'b100011010_000: ratio = -(24'b00000100_1011010001100010);
                        12'b100011010_011: ratio = -(24'b00000100_1000111011001000);
                        12'b100011010_110: ratio = -(24'b00000100_0110101101011011);
                        12'b100011011_001: ratio = -(24'b00000100_0100100111101100);
                        12'b100011011_100: ratio = -(24'b00000100_0010101001010001);
                        12'b100011011_111: ratio = -(24'b00000100_0000110001100011);
                        12'b100011100_010: ratio = -(24'b00000011_1111000000000000);
                        12'b100011100_101: ratio = -(24'b00000011_1101010100001011);
                        12'b100011101_000: ratio = -(24'b00000011_1011101101100111);
                        12'b100011101_011: ratio = -(24'b00000011_1010001011111101);
                        12'b100011101_110: ratio = -(24'b00000011_1000101110110101);
                        12'b100011110_001: ratio = -(24'b00000011_0111010101111011);
                        12'b100011110_100: ratio = -(24'b00000011_0110000000111101);
                        12'b100011110_111: ratio = -(24'b00000011_0100101111101011);
                        12'b100011111_010: ratio = -(24'b00000011_0011100001110100);
                        12'b100011111_101: ratio = -(24'b00000011_0010010111001011);
                        12'b100100000_000: ratio = -(24'b00000011_0001001111100011);
                        12'b100100000_011: ratio = -(24'b00000011_0000001010101111);
                        12'b100100000_110: ratio = -(24'b00000010_1111001000100110);
                        12'b100100001_001: ratio = -(24'b00000010_1110001000111101);
                        12'b100100001_100: ratio = -(24'b00000010_1101001011101011);
                        12'b100100001_111: ratio = -(24'b00000010_1100010000101000);
                        12'b100100010_010: ratio = -(24'b00000010_1011010111101011);
                        12'b100100010_101: ratio = -(24'b00000010_1010100000101100);
                        12'b100100011_000: ratio = -(24'b00000010_1001101011100111);
                        12'b100100011_011: ratio = -(24'b00000010_1000111000010011);
                        12'b100100011_110: ratio = -(24'b00000010_1000000110101011);
                        12'b100100100_001: ratio = -(24'b00000010_0111010110101001);
                        12'b100100100_100: ratio = -(24'b00000010_0110101000001001);
                        12'b100100100_111: ratio = -(24'b00000010_0101111011000110);
                        12'b100100101_010: ratio = -(24'b00000010_0101001111011011);
                        12'b100100101_101: ratio = -(24'b00000010_0100100101000011);
                        12'b100100110_000: ratio = -(24'b00000010_0011111011111100);
                        12'b100100110_011: ratio = -(24'b00000010_0011010100000001);
                        12'b100100110_110: ratio = -(24'b00000010_0010101101001110);
                        12'b100100111_001: ratio = -(24'b00000010_0010000111100001);
                        12'b100100111_100: ratio = -(24'b00000010_0001100010110111);
                        12'b100100111_111: ratio = -(24'b00000010_0000111111001100);
                        12'b100101000_010: ratio = -(24'b00000010_0000011100011101);
                        12'b100101000_101: ratio = -(24'b00000001_1111111010101001);
                        12'b100101001_000: ratio = -(24'b00000001_1111011001101101);
                        12'b100101001_011: ratio = -(24'b00000001_1110111001100110);
                        12'b100101001_110: ratio = -(24'b00000001_1110011010010011);
                        12'b100101010_001: ratio = -(24'b00000001_1101111011110001);
                        12'b100101010_100: ratio = -(24'b00000001_1101011101111110);
                        12'b100101010_111: ratio = -(24'b00000001_1101000000111000);
                        12'b100101011_010: ratio = -(24'b00000001_1100100100011110);
                        12'b100101011_101: ratio = -(24'b00000001_1100001000101111);
                        12'b100101100_000: ratio = -(24'b00000001_1011101101100111);
                        12'b100101100_011: ratio = -(24'b00000001_1011010011000111);
                        12'b100101100_110: ratio = -(24'b00000001_1010111001001100);
                        12'b100101101_001: ratio = -(24'b00000001_1010011111110101);
                        12'b100101101_100: ratio = -(24'b00000001_1010000111000001);
                        12'b100101101_111: ratio = -(24'b00000001_1001101110101110);
                        12'b100101110_010: ratio = -(24'b00000001_1001010110111100);
                        12'b100101110_101: ratio = -(24'b00000001_1000111111101001);
                        12'b100101111_000: ratio = -(24'b00000001_1000101000110100);
                        12'b100101111_011: ratio = -(24'b00000001_1000010010011100);
                        12'b100101111_110: ratio = -(24'b00000001_0111111100100001);
                        12'b100110000_001: ratio = -(24'b00000001_0111100111000001);
                        12'b100110000_100: ratio = -(24'b00000001_0111010001111011);
                        12'b100110000_111: ratio = -(24'b00000001_0110111101001111);
                        12'b100110001_010: ratio = -(24'b00000001_0110101000111011);
                        12'b100110001_101: ratio = -(24'b00000001_0110010100111111);
                        12'b100110010_000: ratio = -(24'b00000001_0110000001011010);
                        12'b100110010_011: ratio = -(24'b00000001_0101101110001100);
                        12'b100110010_110: ratio = -(24'b00000001_0101011011010011);
                        12'b100110011_001: ratio = -(24'b00000001_0101001000101111);
                        12'b100110011_100: ratio = -(24'b00000001_0100110110100000);
                        12'b100110011_111: ratio = -(24'b00000001_0100100100100100);
                        12'b100110100_010: ratio = -(24'b00000001_0100010010111100);
                        12'b100110100_101: ratio = -(24'b00000001_0100000001100110);
                        12'b100110101_000: ratio = -(24'b00000001_0011110000100010);
                        12'b100110101_011: ratio = -(24'b00000001_0011011111101111);
                        12'b100110101_110: ratio = -(24'b00000001_0011001111001110);
                        12'b100110110_001: ratio = -(24'b00000001_0010111110111101);
                        12'b100110110_100: ratio = -(24'b00000001_0010101110111100);
                        12'b100110110_111: ratio = -(24'b00000001_0010011111001011);
                        12'b100110111_010: ratio = -(24'b00000001_0010001111101001);
                        12'b100110111_101: ratio = -(24'b00000001_0010000000010110);
                        12'b100111000_000: ratio = -(24'b00000001_0001110001010001);
                        12'b100111000_011: ratio = -(24'b00000001_0001100010011001);
                        12'b100111000_110: ratio = -(24'b00000001_0001010011110000);
                        12'b100111001_001: ratio = -(24'b00000001_0001000101010100);
                        12'b100111001_100: ratio = -(24'b00000001_0000110111000100);
                        12'b100111001_111: ratio = -(24'b00000001_0000101001000001);
                        12'b100111010_010: ratio = -(24'b00000001_0000011011001010);
                        12'b100111010_101: ratio = -(24'b00000001_0000001101011111);
                        12'b100111011_000: ratio = -(24'b00000000_1111111111111111);
                        12'b100111011_011: ratio = -(24'b00000000_1111110010101011);
                        12'b100111011_110: ratio = -(24'b00000000_1111100101100010);
                        12'b100111100_001: ratio = -(24'b00000000_1111011000100011);
                        12'b100111100_100: ratio = -(24'b00000000_1111001011101111);
                        12'b100111100_111: ratio = -(24'b00000000_1110111111000101);
                        12'b100111101_010: ratio = -(24'b00000000_1110110010100100);
                        12'b100111101_101: ratio = -(24'b00000000_1110100110001110);
                        12'b100111110_000: ratio = -(24'b00000000_1110011010000000);
                        12'b100111110_011: ratio = -(24'b00000000_1110001101111100);
                        12'b100111110_110: ratio = -(24'b00000000_1110000010000001);
                        12'b100111111_001: ratio = -(24'b00000000_1101110110001111);
                        12'b100111111_100: ratio = -(24'b00000000_1101101010100101);
                        12'b100111111_111: ratio = -(24'b00000000_1101011111000011);
                        12'b101000000_010: ratio = -(24'b00000000_1101010011101001);
                        12'b101000000_101: ratio = -(24'b00000000_1101001000011000);
                        12'b101000001_000: ratio = -(24'b00000000_1100111101001110);
                        12'b101000001_011: ratio = -(24'b00000000_1100110010001011);
                        12'b101000001_110: ratio = -(24'b00000000_1100100111010000);
                        12'b101000010_001: ratio = -(24'b00000000_1100011100011100);
                        12'b101000010_100: ratio = -(24'b00000000_1100010001101111);
                        12'b101000010_111: ratio = -(24'b00000000_1100000111001001);
                        12'b101000011_010: ratio = -(24'b00000000_1011111100101010);
                        12'b101000011_101: ratio = -(24'b00000000_1011110010010001);
                        12'b101000100_000: ratio = -(24'b00000000_1011100111111110);
                        12'b101000100_011: ratio = -(24'b00000000_1011011101110010);
                        12'b101000100_110: ratio = -(24'b00000000_1011010011101100);
                        12'b101000101_001: ratio = -(24'b00000000_1011001001101100);
                        12'b101000101_100: ratio = -(24'b00000000_1010111111110001);
                        12'b101000101_111: ratio = -(24'b00000000_1010110101111100);
                        12'b101000110_010: ratio = -(24'b00000000_1010101100001101);
                        12'b101000110_101: ratio = -(24'b00000000_1010100010100100);
                        12'b101000111_000: ratio = -(24'b00000000_1010011000111111);
                        12'b101000111_011: ratio = -(24'b00000000_1010001111100000);
                        12'b101000111_110: ratio = -(24'b00000000_1010000110000110);
                        12'b101001000_001: ratio = -(24'b00000000_1001111100110000);
                        12'b101001000_100: ratio = -(24'b00000000_1001110011100000);
                        12'b101001000_111: ratio = -(24'b00000000_1001101010010100);
                        12'b101001001_010: ratio = -(24'b00000000_1001100001001101);
                        12'b101001001_101: ratio = -(24'b00000000_1001011000001011);
                        12'b101001010_000: ratio = -(24'b00000000_1001001111001101);
                        12'b101001010_011: ratio = -(24'b00000000_1001000110010011);
                        12'b101001010_110: ratio = -(24'b00000000_1000111101011101);
                        12'b101001011_001: ratio = -(24'b00000000_1000110100101100);
                        12'b101001011_100: ratio = -(24'b00000000_1000101011111111);
                        12'b101001011_111: ratio = -(24'b00000000_1000100011010101);
                        12'b101001100_010: ratio = -(24'b00000000_1000011010110000);
                        12'b101001100_101: ratio = -(24'b00000000_1000010010001110);
                        12'b101001101_000: ratio = -(24'b00000000_1000001001110000);
                        12'b101001101_011: ratio = -(24'b00000000_1000000001010101);
                        12'b101001101_110: ratio = -(24'b00000000_0111111000111110);
                        12'b101001110_001: ratio = -(24'b00000000_0111110000101011);
                        12'b101001110_100: ratio = -(24'b00000000_0111101000011011);
                        12'b101001110_111: ratio = -(24'b00000000_0111100000001110);
                        12'b101001111_010: ratio = -(24'b00000000_0111011000000100);
                        12'b101001111_101: ratio = -(24'b00000000_0111001111111101);
                        12'b101010000_000: ratio = -(24'b00000000_0111000111111010);
                        12'b101010000_011: ratio = -(24'b00000000_0110111111111010);
                        12'b101010000_110: ratio = -(24'b00000000_0110110111111100);
                        12'b101010001_001: ratio = -(24'b00000000_0110110000000001);
                        12'b101010001_100: ratio = -(24'b00000000_0110101000001001);
                        12'b101010001_111: ratio = -(24'b00000000_0110100000010100);
                        12'b101010010_010: ratio = -(24'b00000000_0110011000100010);
                        12'b101010010_101: ratio = -(24'b00000000_0110010000110010);
                        12'b101010011_000: ratio = -(24'b00000000_0110001001000100);
                        12'b101010011_011: ratio = -(24'b00000000_0110000001011010);
                        12'b101010011_110: ratio = -(24'b00000000_0101111001110001);
                        12'b101010100_001: ratio = -(24'b00000000_0101110010001011);
                        12'b101010100_100: ratio = -(24'b00000000_0101101010100111);
                        12'b101010100_111: ratio = -(24'b00000000_0101100011000101);
                        12'b101010101_010: ratio = -(24'b00000000_0101011011100110);
                        12'b101010101_101: ratio = -(24'b00000000_0101010100001001);
                        12'b101010110_000: ratio = -(24'b00000000_0101001100101101);
                        12'b101010110_011: ratio = -(24'b00000000_0101000101010100);
                        12'b101010110_110: ratio = -(24'b00000000_0100111101111101);
                        12'b101010111_001: ratio = -(24'b00000000_0100110110101000);
                        12'b101010111_100: ratio = -(24'b00000000_0100101111010100);
                        12'b101010111_111: ratio = -(24'b00000000_0100101000000010);
                        12'b101011000_010: ratio = -(24'b00000000_0100100000110011);
                        12'b101011000_101: ratio = -(24'b00000000_0100011001100100);
                        12'b101011001_000: ratio = -(24'b00000000_0100010010011000);
                        12'b101011001_011: ratio = -(24'b00000000_0100001011001101);
                        12'b101011001_110: ratio = -(24'b00000000_0100000100000100);
                        12'b101011010_001: ratio = -(24'b00000000_0011111100111100);
                        12'b101011010_100: ratio = -(24'b00000000_0011110101110101);
                        12'b101011010_111: ratio = -(24'b00000000_0011101110110000);
                        12'b101011011_010: ratio = -(24'b00000000_0011100111101101);
                        12'b101011011_101: ratio = -(24'b00000000_0011100000101011);
                        12'b101011100_000: ratio = -(24'b00000000_0011011001101010);
                        12'b101011100_011: ratio = -(24'b00000000_0011010010101010);
                        12'b101011100_110: ratio = -(24'b00000000_0011001011101011);
                        12'b101011101_001: ratio = -(24'b00000000_0011000100101110);
                        12'b101011101_100: ratio = -(24'b00000000_0010111101110010);
                        12'b101011101_111: ratio = -(24'b00000000_0010110110110111);
                        12'b101011110_010: ratio = -(24'b00000000_0010101111111101);
                        12'b101011110_101: ratio = -(24'b00000000_0010101001000100);
                        12'b101011111_000: ratio = -(24'b00000000_0010100010001011);
                        12'b101011111_011: ratio = -(24'b00000000_0010011011010100);
                        12'b101011111_110: ratio = -(24'b00000000_0010010100011110);
                        12'b101100000_001: ratio = -(24'b00000000_0010001101101000);
                        12'b101100000_100: ratio = -(24'b00000000_0010000110110011);
                        12'b101100000_111: ratio = -(24'b00000000_0001111111111111);
                        12'b101100001_010: ratio = -(24'b00000000_0001111001001100);
                        12'b101100001_101: ratio = -(24'b00000000_0001110010011010);
                        12'b101100010_000: ratio = -(24'b00000000_0001101011101000);
                        12'b101100010_011: ratio = -(24'b00000000_0001100100110110);
                        12'b101100010_110: ratio = -(24'b00000000_0001011110000101);
                        12'b101100011_001: ratio = -(24'b00000000_0001010111010101);
                        12'b101100011_100: ratio = -(24'b00000000_0001010000100101);
                        12'b101100011_111: ratio = -(24'b00000000_0001001001110110);
                        12'b101100100_010: ratio = -(24'b00000000_0001000011000111);
                        12'b101100100_101: ratio = -(24'b00000000_0000111100011000);
                        12'b101100101_000: ratio = -(24'b00000000_0000110101101010);
                        12'b101100101_011: ratio = -(24'b00000000_0000101110111100);
                        12'b101100101_110: ratio = -(24'b00000000_0000101000001110);
                        12'b101100110_001: ratio = -(24'b00000000_0000100001100001);
                        12'b101100110_100: ratio = -(24'b00000000_0000011010110100);
                        12'b101100110_111: ratio = -(24'b00000000_0000010100000110);
                        12'b101100111_010: ratio = -(24'b00000000_0000001101011001);
                        12'b101100111_101: ratio = -(24'b00000000_0000000110101100);
                        default: ratio = 24'b0;
                endcase
        end
endmodule


