`timescale 1ns/1ns

module raycast_3d_maze(input [3:0] KEY, input [9:0] SW, output [9:0] LEDR);

endmodule
