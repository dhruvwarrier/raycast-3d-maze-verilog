module sin_LUT(input [11:0] angle, output reg [23:0] ratio);

        always @(*) begin
                case(angle)
                        12'b000000000_000: ratio = 24'b00000000_0000000000000000;
                        12'b000000000_011: ratio = 24'b00000000_0000000110101100;
                        12'b000000000_110: ratio = 24'b00000000_0000001101011001;
                        12'b000000001_001: ratio = 24'b00000000_0000010100000110;
                        12'b000000001_100: ratio = 24'b00000000_0000011010110011;
                        12'b000000001_111: ratio = 24'b00000000_0000100001100000;
                        12'b000000010_010: ratio = 24'b00000000_0000101000001100;
                        12'b000000010_101: ratio = 24'b00000000_0000101110111001;
                        12'b000000011_000: ratio = 24'b00000000_0000110101100101;
                        12'b000000011_011: ratio = 24'b00000000_0000111100010010;
                        12'b000000011_110: ratio = 24'b00000000_0001000010111110;
                        12'b000000100_001: ratio = 24'b00000000_0001001001101010;
                        12'b000000100_100: ratio = 24'b00000000_0001010000010101;
                        12'b000000100_111: ratio = 24'b00000000_0001010111000001;
                        12'b000000101_010: ratio = 24'b00000000_0001011101101100;
                        12'b000000101_101: ratio = 24'b00000000_0001100100010111;
                        12'b000000110_000: ratio = 24'b00000000_0001101011000010;
                        12'b000000110_011: ratio = 24'b00000000_0001110001101100;
                        12'b000000110_110: ratio = 24'b00000000_0001111000010110;
                        12'b000000111_001: ratio = 24'b00000000_0001111111000000;
                        12'b000000111_100: ratio = 24'b00000000_0010000101101010;
                        12'b000000111_111: ratio = 24'b00000000_0010001100010011;
                        12'b000001000_010: ratio = 24'b00000000_0010010010111011;
                        12'b000001000_101: ratio = 24'b00000000_0010011001100100;
                        12'b000001001_000: ratio = 24'b00000000_0010100000001100;
                        12'b000001001_011: ratio = 24'b00000000_0010100110110011;
                        12'b000001001_110: ratio = 24'b00000000_0010101101011010;
                        12'b000001010_001: ratio = 24'b00000000_0010110100000000;
                        12'b000001010_100: ratio = 24'b00000000_0010111010100110;
                        12'b000001010_111: ratio = 24'b00000000_0011000001001100;
                        12'b000001011_010: ratio = 24'b00000000_0011000111110001;
                        12'b000001011_101: ratio = 24'b00000000_0011001110010101;
                        12'b000001100_000: ratio = 24'b00000000_0011010100111001;
                        12'b000001100_011: ratio = 24'b00000000_0011011011011100;
                        12'b000001100_110: ratio = 24'b00000000_0011100001111111;
                        12'b000001101_001: ratio = 24'b00000000_0011101000100001;
                        12'b000001101_100: ratio = 24'b00000000_0011101111000011;
                        12'b000001101_111: ratio = 24'b00000000_0011110101100011;
                        12'b000001110_010: ratio = 24'b00000000_0011111100000011;
                        12'b000001110_101: ratio = 24'b00000000_0100000010100011;
                        12'b000001111_000: ratio = 24'b00000000_0100001001000001;
                        12'b000001111_011: ratio = 24'b00000000_0100001111011111;
                        12'b000001111_110: ratio = 24'b00000000_0100010101111101;
                        12'b000010000_001: ratio = 24'b00000000_0100011100011001;
                        12'b000010000_100: ratio = 24'b00000000_0100100010110101;
                        12'b000010000_111: ratio = 24'b00000000_0100101001010000;
                        12'b000010001_010: ratio = 24'b00000000_0100101111101010;
                        12'b000010001_101: ratio = 24'b00000000_0100110110000011;
                        12'b000010010_000: ratio = 24'b00000000_0100111100011011;
                        12'b000010010_011: ratio = 24'b00000000_0101000010110011;
                        12'b000010010_110: ratio = 24'b00000000_0101001001001001;
                        12'b000010011_001: ratio = 24'b00000000_0101001111011111;
                        12'b000010011_100: ratio = 24'b00000000_0101010101110100;
                        12'b000010011_111: ratio = 24'b00000000_0101011100001000;
                        12'b000010100_010: ratio = 24'b00000000_0101100010011011;
                        12'b000010100_101: ratio = 24'b00000000_0101101000101101;
                        12'b000010101_000: ratio = 24'b00000000_0101101110111110;
                        12'b000010101_011: ratio = 24'b00000000_0101110101001101;
                        12'b000010101_110: ratio = 24'b00000000_0101111011011100;
                        12'b000010110_001: ratio = 24'b00000000_0110000001101010;
                        12'b000010110_100: ratio = 24'b00000000_0110000111110111;
                        12'b000010110_111: ratio = 24'b00000000_0110001110000011;
                        12'b000010111_010: ratio = 24'b00000000_0110010100001101;
                        12'b000010111_101: ratio = 24'b00000000_0110011010010111;
                        12'b000011000_000: ratio = 24'b00000000_0110100000011111;
                        12'b000011000_011: ratio = 24'b00000000_0110100110100111;
                        12'b000011000_110: ratio = 24'b00000000_0110101100101101;
                        12'b000011001_001: ratio = 24'b00000000_0110110010110010;
                        12'b000011001_100: ratio = 24'b00000000_0110111000110101;
                        12'b000011001_111: ratio = 24'b00000000_0110111110111000;
                        12'b000011010_010: ratio = 24'b00000000_0111000100111001;
                        12'b000011010_101: ratio = 24'b00000000_0111001010111001;
                        12'b000011011_000: ratio = 24'b00000000_0111010000111000;
                        12'b000011011_011: ratio = 24'b00000000_0111010110110110;
                        12'b000011011_110: ratio = 24'b00000000_0111011100110010;
                        12'b000011100_001: ratio = 24'b00000000_0111100010101101;
                        12'b000011100_100: ratio = 24'b00000000_0111101000100111;
                        12'b000011100_111: ratio = 24'b00000000_0111101110011111;
                        12'b000011101_010: ratio = 24'b00000000_0111110100010110;
                        12'b000011101_101: ratio = 24'b00000000_0111111010001011;
                        12'b000011110_000: ratio = 24'b00000000_1000000000000000;
                        12'b000011110_011: ratio = 24'b00000000_1000000101110010;
                        12'b000011110_110: ratio = 24'b00000000_1000001011100100;
                        12'b000011111_001: ratio = 24'b00000000_1000010001010100;
                        12'b000011111_100: ratio = 24'b00000000_1000010111000010;
                        12'b000011111_111: ratio = 24'b00000000_1000011100101111;
                        12'b000100000_010: ratio = 24'b00000000_1000100010011010;
                        12'b000100000_101: ratio = 24'b00000000_1000101000000100;
                        12'b000100001_000: ratio = 24'b00000000_1000101101101101;
                        12'b000100001_011: ratio = 24'b00000000_1000110011010100;
                        12'b000100001_110: ratio = 24'b00000000_1000111000111001;
                        12'b000100010_001: ratio = 24'b00000000_1000111110011101;
                        12'b000100010_100: ratio = 24'b00000000_1001000011111111;
                        12'b000100010_111: ratio = 24'b00000000_1001001001100000;
                        12'b000100011_010: ratio = 24'b00000000_1001001110111111;
                        12'b000100011_101: ratio = 24'b00000000_1001010100011101;
                        12'b000100100_000: ratio = 24'b00000000_1001011001111001;
                        12'b000100100_011: ratio = 24'b00000000_1001011111010011;
                        12'b000100100_110: ratio = 24'b00000000_1001100100101011;
                        12'b000100101_001: ratio = 24'b00000000_1001101010000010;
                        12'b000100101_100: ratio = 24'b00000000_1001101111010111;
                        12'b000100101_111: ratio = 24'b00000000_1001110100101011;
                        12'b000100110_010: ratio = 24'b00000000_1001111001111100;
                        12'b000100110_101: ratio = 24'b00000000_1001111111001100;
                        12'b000100111_000: ratio = 24'b00000000_1010000100011011;
                        12'b000100111_011: ratio = 24'b00000000_1010001001100111;
                        12'b000100111_110: ratio = 24'b00000000_1010001110110010;
                        12'b000101000_001: ratio = 24'b00000000_1010010011111011;
                        12'b000101000_100: ratio = 24'b00000000_1010011001000010;
                        12'b000101000_111: ratio = 24'b00000000_1010011110000111;
                        12'b000101001_010: ratio = 24'b00000000_1010100011001010;
                        12'b000101001_101: ratio = 24'b00000000_1010101000001100;
                        12'b000101010_000: ratio = 24'b00000000_1010101101001100;
                        12'b000101010_011: ratio = 24'b00000000_1010110010001001;
                        12'b000101010_110: ratio = 24'b00000000_1010110111000101;
                        12'b000101011_001: ratio = 24'b00000000_1010111011111111;
                        12'b000101011_100: ratio = 24'b00000000_1011000000111000;
                        12'b000101011_111: ratio = 24'b00000000_1011000101101110;
                        12'b000101100_010: ratio = 24'b00000000_1011001010100010;
                        12'b000101100_101: ratio = 24'b00000000_1011001111010100;
                        12'b000101101_000: ratio = 24'b00000000_1011010100000100;
                        12'b000101101_011: ratio = 24'b00000000_1011011000110011;
                        12'b000101101_110: ratio = 24'b00000000_1011011101011111;
                        12'b000101110_001: ratio = 24'b00000000_1011100010001001;
                        12'b000101110_100: ratio = 24'b00000000_1011100110110010;
                        12'b000101110_111: ratio = 24'b00000000_1011101011011000;
                        12'b000101111_010: ratio = 24'b00000000_1011101111111100;
                        12'b000101111_101: ratio = 24'b00000000_1011110100011110;
                        12'b000110000_000: ratio = 24'b00000000_1011111000111110;
                        12'b000110000_011: ratio = 24'b00000000_1011111101011100;
                        12'b000110000_110: ratio = 24'b00000000_1100000001111000;
                        12'b000110001_001: ratio = 24'b00000000_1100000110010010;
                        12'b000110001_100: ratio = 24'b00000000_1100001010101001;
                        12'b000110001_111: ratio = 24'b00000000_1100001110111111;
                        12'b000110010_010: ratio = 24'b00000000_1100010011010010;
                        12'b000110010_101: ratio = 24'b00000000_1100010111100100;
                        12'b000110011_000: ratio = 24'b00000000_1100011011110011;
                        12'b000110011_011: ratio = 24'b00000000_1100011111111111;
                        12'b000110011_110: ratio = 24'b00000000_1100100100001010;
                        12'b000110100_001: ratio = 24'b00000000_1100101000010010;
                        12'b000110100_100: ratio = 24'b00000000_1100101100011001;
                        12'b000110100_111: ratio = 24'b00000000_1100110000011101;
                        12'b000110101_010: ratio = 24'b00000000_1100110100011110;
                        12'b000110101_101: ratio = 24'b00000000_1100111000011110;
                        12'b000110110_000: ratio = 24'b00000000_1100111100011011;
                        12'b000110110_011: ratio = 24'b00000000_1101000000010110;
                        12'b000110110_110: ratio = 24'b00000000_1101000100001111;
                        12'b000110111_001: ratio = 24'b00000000_1101001000000101;
                        12'b000110111_100: ratio = 24'b00000000_1101001011111001;
                        12'b000110111_111: ratio = 24'b00000000_1101001111101011;
                        12'b000111000_010: ratio = 24'b00000000_1101010011011011;
                        12'b000111000_101: ratio = 24'b00000000_1101010111001000;
                        12'b000111001_000: ratio = 24'b00000000_1101011010110011;
                        12'b000111001_011: ratio = 24'b00000000_1101011110011011;
                        12'b000111001_110: ratio = 24'b00000000_1101100010000001;
                        12'b000111010_001: ratio = 24'b00000000_1101100101100101;
                        12'b000111010_100: ratio = 24'b00000000_1101101001000110;
                        12'b000111010_111: ratio = 24'b00000000_1101101100100101;
                        12'b000111011_010: ratio = 24'b00000000_1101110000000010;
                        12'b000111011_101: ratio = 24'b00000000_1101110011011100;
                        12'b000111100_000: ratio = 24'b00000000_1101110110110011;
                        12'b000111100_011: ratio = 24'b00000000_1101111010001001;
                        12'b000111100_110: ratio = 24'b00000000_1101111101011011;
                        12'b000111101_001: ratio = 24'b00000000_1110000000101100;
                        12'b000111101_100: ratio = 24'b00000000_1110000011111010;
                        12'b000111101_111: ratio = 24'b00000000_1110000111000101;
                        12'b000111110_010: ratio = 24'b00000000_1110001010001110;
                        12'b000111110_101: ratio = 24'b00000000_1110001101010101;
                        12'b000111111_000: ratio = 24'b00000000_1110010000011001;
                        12'b000111111_011: ratio = 24'b00000000_1110010011011010;
                        12'b000111111_110: ratio = 24'b00000000_1110010110011001;
                        12'b001000000_001: ratio = 24'b00000000_1110011001010101;
                        12'b001000000_100: ratio = 24'b00000000_1110011100001111;
                        12'b001000000_111: ratio = 24'b00000000_1110011111000111;
                        12'b001000001_010: ratio = 24'b00000000_1110100001111100;
                        12'b001000001_101: ratio = 24'b00000000_1110100100101110;
                        12'b001000010_000: ratio = 24'b00000000_1110100111011110;
                        12'b001000010_011: ratio = 24'b00000000_1110101010001011;
                        12'b001000010_110: ratio = 24'b00000000_1110101100110101;
                        12'b001000011_001: ratio = 24'b00000000_1110101111011101;
                        12'b001000011_100: ratio = 24'b00000000_1110110010000011;
                        12'b001000011_111: ratio = 24'b00000000_1110110100100110;
                        12'b001000100_010: ratio = 24'b00000000_1110110111000110;
                        12'b001000100_101: ratio = 24'b00000000_1110111001100100;
                        12'b001000101_000: ratio = 24'b00000000_1110111011111111;
                        12'b001000101_011: ratio = 24'b00000000_1110111110010111;
                        12'b001000101_110: ratio = 24'b00000000_1111000000101101;
                        12'b001000110_001: ratio = 24'b00000000_1111000011000000;
                        12'b001000110_100: ratio = 24'b00000000_1111000101010000;
                        12'b001000110_111: ratio = 24'b00000000_1111000111011110;
                        12'b001000111_010: ratio = 24'b00000000_1111001001101010;
                        12'b001000111_101: ratio = 24'b00000000_1111001011110010;
                        12'b001001000_000: ratio = 24'b00000000_1111001101111000;
                        12'b001001000_011: ratio = 24'b00000000_1111001111111011;
                        12'b001001000_110: ratio = 24'b00000000_1111010001111100;
                        12'b001001001_001: ratio = 24'b00000000_1111010011111010;
                        12'b001001001_100: ratio = 24'b00000000_1111010101110101;
                        12'b001001001_111: ratio = 24'b00000000_1111010111101101;
                        12'b001001010_010: ratio = 24'b00000000_1111011001100011;
                        12'b001001010_101: ratio = 24'b00000000_1111011011010110;
                        12'b001001011_000: ratio = 24'b00000000_1111011101000110;
                        12'b001001011_011: ratio = 24'b00000000_1111011110110100;
                        12'b001001011_110: ratio = 24'b00000000_1111100000011111;
                        12'b001001100_001: ratio = 24'b00000000_1111100010000111;
                        12'b001001100_100: ratio = 24'b00000000_1111100011101101;
                        12'b001001100_111: ratio = 24'b00000000_1111100101010000;
                        12'b001001101_010: ratio = 24'b00000000_1111100110110000;
                        12'b001001101_101: ratio = 24'b00000000_1111101000001101;
                        12'b001001110_000: ratio = 24'b00000000_1111101001100111;
                        12'b001001110_011: ratio = 24'b00000000_1111101010111111;
                        12'b001001110_110: ratio = 24'b00000000_1111101100010100;
                        12'b001001111_001: ratio = 24'b00000000_1111101101100111;
                        12'b001001111_100: ratio = 24'b00000000_1111101110110110;
                        12'b001001111_111: ratio = 24'b00000000_1111110000000011;
                        12'b001010000_010: ratio = 24'b00000000_1111110001001101;
                        12'b001010000_101: ratio = 24'b00000000_1111110010010100;
                        12'b001010001_000: ratio = 24'b00000000_1111110011011001;
                        12'b001010001_011: ratio = 24'b00000000_1111110100011010;
                        12'b001010001_110: ratio = 24'b00000000_1111110101011001;
                        12'b001010010_001: ratio = 24'b00000000_1111110110010101;
                        12'b001010010_100: ratio = 24'b00000000_1111110111001111;
                        12'b001010010_111: ratio = 24'b00000000_1111111000000101;
                        12'b001010011_010: ratio = 24'b00000000_1111111000111001;
                        12'b001010011_101: ratio = 24'b00000000_1111111001101010;
                        12'b001010100_000: ratio = 24'b00000000_1111111010011000;
                        12'b001010100_011: ratio = 24'b00000000_1111111011000100;
                        12'b001010100_110: ratio = 24'b00000000_1111111011101101;
                        12'b001010101_001: ratio = 24'b00000000_1111111100010010;
                        12'b001010101_100: ratio = 24'b00000000_1111111100110101;
                        12'b001010101_111: ratio = 24'b00000000_1111111101010110;
                        12'b001010110_010: ratio = 24'b00000000_1111111101110011;
                        12'b001010110_101: ratio = 24'b00000000_1111111110001110;
                        12'b001010111_000: ratio = 24'b00000000_1111111110100110;
                        12'b001010111_011: ratio = 24'b00000000_1111111110111011;
                        12'b001010111_110: ratio = 24'b00000000_1111111111001101;
                        12'b001011000_001: ratio = 24'b00000000_1111111111011100;
                        12'b001011000_100: ratio = 24'b00000000_1111111111101001;
                        12'b001011000_111: ratio = 24'b00000000_1111111111110011;
                        12'b001011001_010: ratio = 24'b00000000_1111111111111010;
                        12'b001011001_101: ratio = 24'b00000000_1111111111111110;
                        12'b001011010_000: ratio = 24'b00000001_0000000000000000;
                        12'b001011010_011: ratio = 24'b00000000_1111111111111110;
                        12'b001011010_110: ratio = 24'b00000000_1111111111111010;
                        12'b001011011_001: ratio = 24'b00000000_1111111111110011;
                        12'b001011011_100: ratio = 24'b00000000_1111111111101001;
                        12'b001011011_111: ratio = 24'b00000000_1111111111011100;
                        12'b001011100_010: ratio = 24'b00000000_1111111111001101;
                        12'b001011100_101: ratio = 24'b00000000_1111111110111011;
                        12'b001011101_000: ratio = 24'b00000000_1111111110100110;
                        12'b001011101_011: ratio = 24'b00000000_1111111110001110;
                        12'b001011101_110: ratio = 24'b00000000_1111111101110011;
                        12'b001011110_001: ratio = 24'b00000000_1111111101010110;
                        12'b001011110_100: ratio = 24'b00000000_1111111100110101;
                        12'b001011110_111: ratio = 24'b00000000_1111111100010010;
                        12'b001011111_010: ratio = 24'b00000000_1111111011101101;
                        12'b001011111_101: ratio = 24'b00000000_1111111011000100;
                        12'b001100000_000: ratio = 24'b00000000_1111111010011000;
                        12'b001100000_011: ratio = 24'b00000000_1111111001101010;
                        12'b001100000_110: ratio = 24'b00000000_1111111000111001;
                        12'b001100001_001: ratio = 24'b00000000_1111111000000101;
                        12'b001100001_100: ratio = 24'b00000000_1111110111001111;
                        12'b001100001_111: ratio = 24'b00000000_1111110110010101;
                        12'b001100010_010: ratio = 24'b00000000_1111110101011001;
                        12'b001100010_101: ratio = 24'b00000000_1111110100011010;
                        12'b001100011_000: ratio = 24'b00000000_1111110011011001;
                        12'b001100011_011: ratio = 24'b00000000_1111110010010100;
                        12'b001100011_110: ratio = 24'b00000000_1111110001001101;
                        12'b001100100_001: ratio = 24'b00000000_1111110000000011;
                        12'b001100100_100: ratio = 24'b00000000_1111101110110110;
                        12'b001100100_111: ratio = 24'b00000000_1111101101100111;
                        12'b001100101_010: ratio = 24'b00000000_1111101100010100;
                        12'b001100101_101: ratio = 24'b00000000_1111101010111111;
                        12'b001100110_000: ratio = 24'b00000000_1111101001100111;
                        12'b001100110_011: ratio = 24'b00000000_1111101000001101;
                        12'b001100110_110: ratio = 24'b00000000_1111100110110000;
                        12'b001100111_001: ratio = 24'b00000000_1111100101010000;
                        12'b001100111_100: ratio = 24'b00000000_1111100011101101;
                        12'b001100111_111: ratio = 24'b00000000_1111100010000111;
                        12'b001101000_010: ratio = 24'b00000000_1111100000011111;
                        12'b001101000_101: ratio = 24'b00000000_1111011110110100;
                        12'b001101001_000: ratio = 24'b00000000_1111011101000110;
                        12'b001101001_011: ratio = 24'b00000000_1111011011010110;
                        12'b001101001_110: ratio = 24'b00000000_1111011001100011;
                        12'b001101010_001: ratio = 24'b00000000_1111010111101101;
                        12'b001101010_100: ratio = 24'b00000000_1111010101110101;
                        12'b001101010_111: ratio = 24'b00000000_1111010011111010;
                        12'b001101011_010: ratio = 24'b00000000_1111010001111100;
                        12'b001101011_101: ratio = 24'b00000000_1111001111111011;
                        12'b001101100_000: ratio = 24'b00000000_1111001101111000;
                        12'b001101100_011: ratio = 24'b00000000_1111001011110010;
                        12'b001101100_110: ratio = 24'b00000000_1111001001101010;
                        12'b001101101_001: ratio = 24'b00000000_1111000111011110;
                        12'b001101101_100: ratio = 24'b00000000_1111000101010000;
                        12'b001101101_111: ratio = 24'b00000000_1111000011000000;
                        12'b001101110_010: ratio = 24'b00000000_1111000000101101;
                        12'b001101110_101: ratio = 24'b00000000_1110111110010111;
                        12'b001101111_000: ratio = 24'b00000000_1110111011111111;
                        12'b001101111_011: ratio = 24'b00000000_1110111001100100;
                        12'b001101111_110: ratio = 24'b00000000_1110110111000110;
                        12'b001110000_001: ratio = 24'b00000000_1110110100100110;
                        12'b001110000_100: ratio = 24'b00000000_1110110010000011;
                        12'b001110000_111: ratio = 24'b00000000_1110101111011101;
                        12'b001110001_010: ratio = 24'b00000000_1110101100110101;
                        12'b001110001_101: ratio = 24'b00000000_1110101010001011;
                        12'b001110010_000: ratio = 24'b00000000_1110100111011110;
                        12'b001110010_011: ratio = 24'b00000000_1110100100101110;
                        12'b001110010_110: ratio = 24'b00000000_1110100001111100;
                        12'b001110011_001: ratio = 24'b00000000_1110011111000111;
                        12'b001110011_100: ratio = 24'b00000000_1110011100001111;
                        12'b001110011_111: ratio = 24'b00000000_1110011001010101;
                        12'b001110100_010: ratio = 24'b00000000_1110010110011001;
                        12'b001110100_101: ratio = 24'b00000000_1110010011011010;
                        12'b001110101_000: ratio = 24'b00000000_1110010000011001;
                        12'b001110101_011: ratio = 24'b00000000_1110001101010101;
                        12'b001110101_110: ratio = 24'b00000000_1110001010001110;
                        12'b001110110_001: ratio = 24'b00000000_1110000111000101;
                        12'b001110110_100: ratio = 24'b00000000_1110000011111010;
                        12'b001110110_111: ratio = 24'b00000000_1110000000101100;
                        12'b001110111_010: ratio = 24'b00000000_1101111101011011;
                        12'b001110111_101: ratio = 24'b00000000_1101111010001001;
                        12'b001111000_000: ratio = 24'b00000000_1101110110110011;
                        12'b001111000_011: ratio = 24'b00000000_1101110011011100;
                        12'b001111000_110: ratio = 24'b00000000_1101110000000010;
                        12'b001111001_001: ratio = 24'b00000000_1101101100100101;
                        12'b001111001_100: ratio = 24'b00000000_1101101001000110;
                        12'b001111001_111: ratio = 24'b00000000_1101100101100101;
                        12'b001111010_010: ratio = 24'b00000000_1101100010000001;
                        12'b001111010_101: ratio = 24'b00000000_1101011110011011;
                        12'b001111011_000: ratio = 24'b00000000_1101011010110011;
                        12'b001111011_011: ratio = 24'b00000000_1101010111001000;
                        12'b001111011_110: ratio = 24'b00000000_1101010011011011;
                        12'b001111100_001: ratio = 24'b00000000_1101001111101011;
                        12'b001111100_100: ratio = 24'b00000000_1101001011111001;
                        12'b001111100_111: ratio = 24'b00000000_1101001000000101;
                        12'b001111101_010: ratio = 24'b00000000_1101000100001111;
                        12'b001111101_101: ratio = 24'b00000000_1101000000010110;
                        12'b001111110_000: ratio = 24'b00000000_1100111100011011;
                        12'b001111110_011: ratio = 24'b00000000_1100111000011110;
                        12'b001111110_110: ratio = 24'b00000000_1100110100011110;
                        12'b001111111_001: ratio = 24'b00000000_1100110000011101;
                        12'b001111111_100: ratio = 24'b00000000_1100101100011001;
                        12'b001111111_111: ratio = 24'b00000000_1100101000010010;
                        12'b010000000_010: ratio = 24'b00000000_1100100100001010;
                        12'b010000000_101: ratio = 24'b00000000_1100011111111111;
                        12'b010000001_000: ratio = 24'b00000000_1100011011110011;
                        12'b010000001_011: ratio = 24'b00000000_1100010111100100;
                        12'b010000001_110: ratio = 24'b00000000_1100010011010010;
                        12'b010000010_001: ratio = 24'b00000000_1100001110111111;
                        12'b010000010_100: ratio = 24'b00000000_1100001010101001;
                        12'b010000010_111: ratio = 24'b00000000_1100000110010010;
                        12'b010000011_010: ratio = 24'b00000000_1100000001111000;
                        12'b010000011_101: ratio = 24'b00000000_1011111101011100;
                        12'b010000100_000: ratio = 24'b00000000_1011111000111110;
                        12'b010000100_011: ratio = 24'b00000000_1011110100011110;
                        12'b010000100_110: ratio = 24'b00000000_1011101111111100;
                        12'b010000101_001: ratio = 24'b00000000_1011101011011000;
                        12'b010000101_100: ratio = 24'b00000000_1011100110110010;
                        12'b010000101_111: ratio = 24'b00000000_1011100010001001;
                        12'b010000110_010: ratio = 24'b00000000_1011011101011111;
                        12'b010000110_101: ratio = 24'b00000000_1011011000110011;
                        12'b010000111_000: ratio = 24'b00000000_1011010100000100;
                        12'b010000111_011: ratio = 24'b00000000_1011001111010100;
                        12'b010000111_110: ratio = 24'b00000000_1011001010100010;
                        12'b010001000_001: ratio = 24'b00000000_1011000101101110;
                        12'b010001000_100: ratio = 24'b00000000_1011000000111000;
                        12'b010001000_111: ratio = 24'b00000000_1010111011111111;
                        12'b010001001_010: ratio = 24'b00000000_1010110111000101;
                        12'b010001001_101: ratio = 24'b00000000_1010110010001001;
                        12'b010001010_000: ratio = 24'b00000000_1010101101001100;
                        12'b010001010_011: ratio = 24'b00000000_1010101000001100;
                        12'b010001010_110: ratio = 24'b00000000_1010100011001010;
                        12'b010001011_001: ratio = 24'b00000000_1010011110000111;
                        12'b010001011_100: ratio = 24'b00000000_1010011001000010;
                        12'b010001011_111: ratio = 24'b00000000_1010010011111011;
                        12'b010001100_010: ratio = 24'b00000000_1010001110110010;
                        12'b010001100_101: ratio = 24'b00000000_1010001001100111;
                        12'b010001101_000: ratio = 24'b00000000_1010000100011011;
                        12'b010001101_011: ratio = 24'b00000000_1001111111001100;
                        12'b010001101_110: ratio = 24'b00000000_1001111001111100;
                        12'b010001110_001: ratio = 24'b00000000_1001110100101011;
                        12'b010001110_100: ratio = 24'b00000000_1001101111010111;
                        12'b010001110_111: ratio = 24'b00000000_1001101010000010;
                        12'b010001111_010: ratio = 24'b00000000_1001100100101011;
                        12'b010001111_101: ratio = 24'b00000000_1001011111010011;
                        12'b010010000_000: ratio = 24'b00000000_1001011001111001;
                        12'b010010000_011: ratio = 24'b00000000_1001010100011101;
                        12'b010010000_110: ratio = 24'b00000000_1001001110111111;
                        12'b010010001_001: ratio = 24'b00000000_1001001001100000;
                        12'b010010001_100: ratio = 24'b00000000_1001000011111111;
                        12'b010010001_111: ratio = 24'b00000000_1000111110011101;
                        12'b010010010_010: ratio = 24'b00000000_1000111000111001;
                        12'b010010010_101: ratio = 24'b00000000_1000110011010100;
                        12'b010010011_000: ratio = 24'b00000000_1000101101101101;
                        12'b010010011_011: ratio = 24'b00000000_1000101000000100;
                        12'b010010011_110: ratio = 24'b00000000_1000100010011010;
                        12'b010010100_001: ratio = 24'b00000000_1000011100101111;
                        12'b010010100_100: ratio = 24'b00000000_1000010111000010;
                        12'b010010100_111: ratio = 24'b00000000_1000010001010100;
                        12'b010010101_010: ratio = 24'b00000000_1000001011100100;
                        12'b010010101_101: ratio = 24'b00000000_1000000101110010;
                        12'b010010110_000: ratio = 24'b00000000_0111111111111111;
                        12'b010010110_011: ratio = 24'b00000000_0111111010001011;
                        12'b010010110_110: ratio = 24'b00000000_0111110100010110;
                        12'b010010111_001: ratio = 24'b00000000_0111101110011111;
                        12'b010010111_100: ratio = 24'b00000000_0111101000100111;
                        12'b010010111_111: ratio = 24'b00000000_0111100010101101;
                        12'b010011000_010: ratio = 24'b00000000_0111011100110010;
                        12'b010011000_101: ratio = 24'b00000000_0111010110110110;
                        12'b010011001_000: ratio = 24'b00000000_0111010000111000;
                        12'b010011001_011: ratio = 24'b00000000_0111001010111001;
                        12'b010011001_110: ratio = 24'b00000000_0111000100111001;
                        12'b010011010_001: ratio = 24'b00000000_0110111110111000;
                        12'b010011010_100: ratio = 24'b00000000_0110111000110101;
                        12'b010011010_111: ratio = 24'b00000000_0110110010110010;
                        12'b010011011_010: ratio = 24'b00000000_0110101100101101;
                        12'b010011011_101: ratio = 24'b00000000_0110100110100111;
                        12'b010011100_000: ratio = 24'b00000000_0110100000011111;
                        12'b010011100_011: ratio = 24'b00000000_0110011010010111;
                        12'b010011100_110: ratio = 24'b00000000_0110010100001101;
                        12'b010011101_001: ratio = 24'b00000000_0110001110000011;
                        12'b010011101_100: ratio = 24'b00000000_0110000111110111;
                        12'b010011101_111: ratio = 24'b00000000_0110000001101010;
                        12'b010011110_010: ratio = 24'b00000000_0101111011011100;
                        12'b010011110_101: ratio = 24'b00000000_0101110101001101;
                        12'b010011111_000: ratio = 24'b00000000_0101101110111110;
                        12'b010011111_011: ratio = 24'b00000000_0101101000101101;
                        12'b010011111_110: ratio = 24'b00000000_0101100010011011;
                        12'b010100000_001: ratio = 24'b00000000_0101011100001000;
                        12'b010100000_100: ratio = 24'b00000000_0101010101110100;
                        12'b010100000_111: ratio = 24'b00000000_0101001111011111;
                        12'b010100001_010: ratio = 24'b00000000_0101001001001001;
                        12'b010100001_101: ratio = 24'b00000000_0101000010110011;
                        12'b010100010_000: ratio = 24'b00000000_0100111100011011;
                        12'b010100010_011: ratio = 24'b00000000_0100110110000011;
                        12'b010100010_110: ratio = 24'b00000000_0100101111101010;
                        12'b010100011_001: ratio = 24'b00000000_0100101001010000;
                        12'b010100011_100: ratio = 24'b00000000_0100100010110101;
                        12'b010100011_111: ratio = 24'b00000000_0100011100011001;
                        12'b010100100_010: ratio = 24'b00000000_0100010101111101;
                        12'b010100100_101: ratio = 24'b00000000_0100001111011111;
                        12'b010100101_000: ratio = 24'b00000000_0100001001000001;
                        12'b010100101_011: ratio = 24'b00000000_0100000010100011;
                        12'b010100101_110: ratio = 24'b00000000_0011111100000011;
                        12'b010100110_001: ratio = 24'b00000000_0011110101100011;
                        12'b010100110_100: ratio = 24'b00000000_0011101111000011;
                        12'b010100110_111: ratio = 24'b00000000_0011101000100001;
                        12'b010100111_010: ratio = 24'b00000000_0011100001111111;
                        12'b010100111_101: ratio = 24'b00000000_0011011011011100;
                        12'b010101000_000: ratio = 24'b00000000_0011010100111001;
                        12'b010101000_011: ratio = 24'b00000000_0011001110010101;
                        12'b010101000_110: ratio = 24'b00000000_0011000111110001;
                        12'b010101001_001: ratio = 24'b00000000_0011000001001100;
                        12'b010101001_100: ratio = 24'b00000000_0010111010100110;
                        12'b010101001_111: ratio = 24'b00000000_0010110100000000;
                        12'b010101010_010: ratio = 24'b00000000_0010101101011010;
                        12'b010101010_101: ratio = 24'b00000000_0010100110110011;
                        12'b010101011_000: ratio = 24'b00000000_0010100000001100;
                        12'b010101011_011: ratio = 24'b00000000_0010011001100100;
                        12'b010101011_110: ratio = 24'b00000000_0010010010111011;
                        12'b010101100_001: ratio = 24'b00000000_0010001100010011;
                        12'b010101100_100: ratio = 24'b00000000_0010000101101010;
                        12'b010101100_111: ratio = 24'b00000000_0001111111000000;
                        12'b010101101_010: ratio = 24'b00000000_0001111000010110;
                        12'b010101101_101: ratio = 24'b00000000_0001110001101100;
                        12'b010101110_000: ratio = 24'b00000000_0001101011000010;
                        12'b010101110_011: ratio = 24'b00000000_0001100100010111;
                        12'b010101110_110: ratio = 24'b00000000_0001011101101100;
                        12'b010101111_001: ratio = 24'b00000000_0001010111000001;
                        12'b010101111_100: ratio = 24'b00000000_0001010000010101;
                        12'b010101111_111: ratio = 24'b00000000_0001001001101010;
                        12'b010110000_010: ratio = 24'b00000000_0001000010111110;
                        12'b010110000_101: ratio = 24'b00000000_0000111100010010;
                        12'b010110001_000: ratio = 24'b00000000_0000110101100101;
                        12'b010110001_011: ratio = 24'b00000000_0000101110111001;
                        12'b010110001_110: ratio = 24'b00000000_0000101000001100;
                        12'b010110010_001: ratio = 24'b00000000_0000100001100000;
                        12'b010110010_100: ratio = 24'b00000000_0000011010110011;
                        12'b010110010_111: ratio = 24'b00000000_0000010100000110;
                        12'b010110011_010: ratio = 24'b00000000_0000001101011001;
                        12'b010110011_101: ratio = 24'b00000000_0000000110101100;
                        12'b010110100_000: ratio = -(24'b00000000_0000000000000000);
                        12'b010110100_011: ratio = -(24'b00000000_0000000110101100);
                        12'b010110100_110: ratio = -(24'b00000000_0000001101011001);
                        12'b010110101_001: ratio = -(24'b00000000_0000010100000110);
                        12'b010110101_100: ratio = -(24'b00000000_0000011010110011);
                        12'b010110101_111: ratio = -(24'b00000000_0000100001100000);
                        12'b010110110_010: ratio = -(24'b00000000_0000101000001100);
                        12'b010110110_101: ratio = -(24'b00000000_0000101110111001);
                        12'b010110111_000: ratio = -(24'b00000000_0000110101100101);
                        12'b010110111_011: ratio = -(24'b00000000_0000111100010010);
                        12'b010110111_110: ratio = -(24'b00000000_0001000010111110);
                        12'b010111000_001: ratio = -(24'b00000000_0001001001101010);
                        12'b010111000_100: ratio = -(24'b00000000_0001010000010101);
                        12'b010111000_111: ratio = -(24'b00000000_0001010111000001);
                        12'b010111001_010: ratio = -(24'b00000000_0001011101101100);
                        12'b010111001_101: ratio = -(24'b00000000_0001100100010111);
                        12'b010111010_000: ratio = -(24'b00000000_0001101011000010);
                        12'b010111010_011: ratio = -(24'b00000000_0001110001101100);
                        12'b010111010_110: ratio = -(24'b00000000_0001111000010110);
                        12'b010111011_001: ratio = -(24'b00000000_0001111111000000);
                        12'b010111011_100: ratio = -(24'b00000000_0010000101101010);
                        12'b010111011_111: ratio = -(24'b00000000_0010001100010011);
                        12'b010111100_010: ratio = -(24'b00000000_0010010010111011);
                        12'b010111100_101: ratio = -(24'b00000000_0010011001100100);
                        12'b010111101_000: ratio = -(24'b00000000_0010100000001100);
                        12'b010111101_011: ratio = -(24'b00000000_0010100110110011);
                        12'b010111101_110: ratio = -(24'b00000000_0010101101011010);
                        12'b010111110_001: ratio = -(24'b00000000_0010110100000000);
                        12'b010111110_100: ratio = -(24'b00000000_0010111010100110);
                        12'b010111110_111: ratio = -(24'b00000000_0011000001001100);
                        12'b010111111_010: ratio = -(24'b00000000_0011000111110001);
                        12'b010111111_101: ratio = -(24'b00000000_0011001110010101);
                        12'b011000000_000: ratio = -(24'b00000000_0011010100111001);
                        12'b011000000_011: ratio = -(24'b00000000_0011011011011100);
                        12'b011000000_110: ratio = -(24'b00000000_0011100001111111);
                        12'b011000001_001: ratio = -(24'b00000000_0011101000100001);
                        12'b011000001_100: ratio = -(24'b00000000_0011101111000011);
                        12'b011000001_111: ratio = -(24'b00000000_0011110101100011);
                        12'b011000010_010: ratio = -(24'b00000000_0011111100000011);
                        12'b011000010_101: ratio = -(24'b00000000_0100000010100011);
                        12'b011000011_000: ratio = -(24'b00000000_0100001001000001);
                        12'b011000011_011: ratio = -(24'b00000000_0100001111011111);
                        12'b011000011_110: ratio = -(24'b00000000_0100010101111101);
                        12'b011000100_001: ratio = -(24'b00000000_0100011100011001);
                        12'b011000100_100: ratio = -(24'b00000000_0100100010110101);
                        12'b011000100_111: ratio = -(24'b00000000_0100101001010000);
                        12'b011000101_010: ratio = -(24'b00000000_0100101111101010);
                        12'b011000101_101: ratio = -(24'b00000000_0100110110000011);
                        12'b011000110_000: ratio = -(24'b00000000_0100111100011011);
                        12'b011000110_011: ratio = -(24'b00000000_0101000010110011);
                        12'b011000110_110: ratio = -(24'b00000000_0101001001001001);
                        12'b011000111_001: ratio = -(24'b00000000_0101001111011111);
                        12'b011000111_100: ratio = -(24'b00000000_0101010101110100);
                        12'b011000111_111: ratio = -(24'b00000000_0101011100001000);
                        12'b011001000_010: ratio = -(24'b00000000_0101100010011011);
                        12'b011001000_101: ratio = -(24'b00000000_0101101000101101);
                        12'b011001001_000: ratio = -(24'b00000000_0101101110111110);
                        12'b011001001_011: ratio = -(24'b00000000_0101110101001101);
                        12'b011001001_110: ratio = -(24'b00000000_0101111011011100);
                        12'b011001010_001: ratio = -(24'b00000000_0110000001101010);
                        12'b011001010_100: ratio = -(24'b00000000_0110000111110111);
                        12'b011001010_111: ratio = -(24'b00000000_0110001110000011);
                        12'b011001011_010: ratio = -(24'b00000000_0110010100001101);
                        12'b011001011_101: ratio = -(24'b00000000_0110011010010111);
                        12'b011001100_000: ratio = -(24'b00000000_0110100000011111);
                        12'b011001100_011: ratio = -(24'b00000000_0110100110100111);
                        12'b011001100_110: ratio = -(24'b00000000_0110101100101101);
                        12'b011001101_001: ratio = -(24'b00000000_0110110010110010);
                        12'b011001101_100: ratio = -(24'b00000000_0110111000110101);
                        12'b011001101_111: ratio = -(24'b00000000_0110111110111000);
                        12'b011001110_010: ratio = -(24'b00000000_0111000100111001);
                        12'b011001110_101: ratio = -(24'b00000000_0111001010111001);
                        12'b011001111_000: ratio = -(24'b00000000_0111010000111000);
                        12'b011001111_011: ratio = -(24'b00000000_0111010110110110);
                        12'b011001111_110: ratio = -(24'b00000000_0111011100110010);
                        12'b011010000_001: ratio = -(24'b00000000_0111100010101101);
                        12'b011010000_100: ratio = -(24'b00000000_0111101000100111);
                        12'b011010000_111: ratio = -(24'b00000000_0111101110011111);
                        12'b011010001_010: ratio = -(24'b00000000_0111110100010110);
                        12'b011010001_101: ratio = -(24'b00000000_0111111010001011);
                        12'b011010010_000: ratio = -(24'b00000000_1000000000000000);
                        12'b011010010_011: ratio = -(24'b00000000_1000000101110010);
                        12'b011010010_110: ratio = -(24'b00000000_1000001011100100);
                        12'b011010011_001: ratio = -(24'b00000000_1000010001010100);
                        12'b011010011_100: ratio = -(24'b00000000_1000010111000010);
                        12'b011010011_111: ratio = -(24'b00000000_1000011100101111);
                        12'b011010100_010: ratio = -(24'b00000000_1000100010011010);
                        12'b011010100_101: ratio = -(24'b00000000_1000101000000100);
                        12'b011010101_000: ratio = -(24'b00000000_1000101101101101);
                        12'b011010101_011: ratio = -(24'b00000000_1000110011010100);
                        12'b011010101_110: ratio = -(24'b00000000_1000111000111001);
                        12'b011010110_001: ratio = -(24'b00000000_1000111110011101);
                        12'b011010110_100: ratio = -(24'b00000000_1001000011111111);
                        12'b011010110_111: ratio = -(24'b00000000_1001001001100000);
                        12'b011010111_010: ratio = -(24'b00000000_1001001110111111);
                        12'b011010111_101: ratio = -(24'b00000000_1001010100011101);
                        12'b011011000_000: ratio = -(24'b00000000_1001011001111001);
                        12'b011011000_011: ratio = -(24'b00000000_1001011111010011);
                        12'b011011000_110: ratio = -(24'b00000000_1001100100101011);
                        12'b011011001_001: ratio = -(24'b00000000_1001101010000010);
                        12'b011011001_100: ratio = -(24'b00000000_1001101111010111);
                        12'b011011001_111: ratio = -(24'b00000000_1001110100101011);
                        12'b011011010_010: ratio = -(24'b00000000_1001111001111100);
                        12'b011011010_101: ratio = -(24'b00000000_1001111111001100);
                        12'b011011011_000: ratio = -(24'b00000000_1010000100011011);
                        12'b011011011_011: ratio = -(24'b00000000_1010001001100111);
                        12'b011011011_110: ratio = -(24'b00000000_1010001110110010);
                        12'b011011100_001: ratio = -(24'b00000000_1010010011111011);
                        12'b011011100_100: ratio = -(24'b00000000_1010011001000010);
                        12'b011011100_111: ratio = -(24'b00000000_1010011110000111);
                        12'b011011101_010: ratio = -(24'b00000000_1010100011001010);
                        12'b011011101_101: ratio = -(24'b00000000_1010101000001100);
                        12'b011011110_000: ratio = -(24'b00000000_1010101101001100);
                        12'b011011110_011: ratio = -(24'b00000000_1010110010001001);
                        12'b011011110_110: ratio = -(24'b00000000_1010110111000101);
                        12'b011011111_001: ratio = -(24'b00000000_1010111011111111);
                        12'b011011111_100: ratio = -(24'b00000000_1011000000111000);
                        12'b011011111_111: ratio = -(24'b00000000_1011000101101110);
                        12'b011100000_010: ratio = -(24'b00000000_1011001010100010);
                        12'b011100000_101: ratio = -(24'b00000000_1011001111010100);
                        12'b011100001_000: ratio = -(24'b00000000_1011010100000100);
                        12'b011100001_011: ratio = -(24'b00000000_1011011000110011);
                        12'b011100001_110: ratio = -(24'b00000000_1011011101011111);
                        12'b011100010_001: ratio = -(24'b00000000_1011100010001001);
                        12'b011100010_100: ratio = -(24'b00000000_1011100110110010);
                        12'b011100010_111: ratio = -(24'b00000000_1011101011011000);
                        12'b011100011_010: ratio = -(24'b00000000_1011101111111100);
                        12'b011100011_101: ratio = -(24'b00000000_1011110100011110);
                        12'b011100100_000: ratio = -(24'b00000000_1011111000111110);
                        12'b011100100_011: ratio = -(24'b00000000_1011111101011100);
                        12'b011100100_110: ratio = -(24'b00000000_1100000001111000);
                        12'b011100101_001: ratio = -(24'b00000000_1100000110010010);
                        12'b011100101_100: ratio = -(24'b00000000_1100001010101001);
                        12'b011100101_111: ratio = -(24'b00000000_1100001110111111);
                        12'b011100110_010: ratio = -(24'b00000000_1100010011010010);
                        12'b011100110_101: ratio = -(24'b00000000_1100010111100100);
                        12'b011100111_000: ratio = -(24'b00000000_1100011011110011);
                        12'b011100111_011: ratio = -(24'b00000000_1100011111111111);
                        12'b011100111_110: ratio = -(24'b00000000_1100100100001010);
                        12'b011101000_001: ratio = -(24'b00000000_1100101000010010);
                        12'b011101000_100: ratio = -(24'b00000000_1100101100011001);
                        12'b011101000_111: ratio = -(24'b00000000_1100110000011101);
                        12'b011101001_010: ratio = -(24'b00000000_1100110100011110);
                        12'b011101001_101: ratio = -(24'b00000000_1100111000011110);
                        12'b011101010_000: ratio = -(24'b00000000_1100111100011011);
                        12'b011101010_011: ratio = -(24'b00000000_1101000000010110);
                        12'b011101010_110: ratio = -(24'b00000000_1101000100001111);
                        12'b011101011_001: ratio = -(24'b00000000_1101001000000101);
                        12'b011101011_100: ratio = -(24'b00000000_1101001011111001);
                        12'b011101011_111: ratio = -(24'b00000000_1101001111101011);
                        12'b011101100_010: ratio = -(24'b00000000_1101010011011011);
                        12'b011101100_101: ratio = -(24'b00000000_1101010111001000);
                        12'b011101101_000: ratio = -(24'b00000000_1101011010110011);
                        12'b011101101_011: ratio = -(24'b00000000_1101011110011011);
                        12'b011101101_110: ratio = -(24'b00000000_1101100010000001);
                        12'b011101110_001: ratio = -(24'b00000000_1101100101100101);
                        12'b011101110_100: ratio = -(24'b00000000_1101101001000110);
                        12'b011101110_111: ratio = -(24'b00000000_1101101100100101);
                        12'b011101111_010: ratio = -(24'b00000000_1101110000000010);
                        12'b011101111_101: ratio = -(24'b00000000_1101110011011100);
                        12'b011110000_000: ratio = -(24'b00000000_1101110110110011);
                        12'b011110000_011: ratio = -(24'b00000000_1101111010001001);
                        12'b011110000_110: ratio = -(24'b00000000_1101111101011011);
                        12'b011110001_001: ratio = -(24'b00000000_1110000000101100);
                        12'b011110001_100: ratio = -(24'b00000000_1110000011111010);
                        12'b011110001_111: ratio = -(24'b00000000_1110000111000101);
                        12'b011110010_010: ratio = -(24'b00000000_1110001010001110);
                        12'b011110010_101: ratio = -(24'b00000000_1110001101010101);
                        12'b011110011_000: ratio = -(24'b00000000_1110010000011001);
                        12'b011110011_011: ratio = -(24'b00000000_1110010011011010);
                        12'b011110011_110: ratio = -(24'b00000000_1110010110011001);
                        12'b011110100_001: ratio = -(24'b00000000_1110011001010101);
                        12'b011110100_100: ratio = -(24'b00000000_1110011100001111);
                        12'b011110100_111: ratio = -(24'b00000000_1110011111000111);
                        12'b011110101_010: ratio = -(24'b00000000_1110100001111100);
                        12'b011110101_101: ratio = -(24'b00000000_1110100100101110);
                        12'b011110110_000: ratio = -(24'b00000000_1110100111011110);
                        12'b011110110_011: ratio = -(24'b00000000_1110101010001011);
                        12'b011110110_110: ratio = -(24'b00000000_1110101100110101);
                        12'b011110111_001: ratio = -(24'b00000000_1110101111011101);
                        12'b011110111_100: ratio = -(24'b00000000_1110110010000011);
                        12'b011110111_111: ratio = -(24'b00000000_1110110100100110);
                        12'b011111000_010: ratio = -(24'b00000000_1110110111000110);
                        12'b011111000_101: ratio = -(24'b00000000_1110111001100100);
                        12'b011111001_000: ratio = -(24'b00000000_1110111011111111);
                        12'b011111001_011: ratio = -(24'b00000000_1110111110010111);
                        12'b011111001_110: ratio = -(24'b00000000_1111000000101101);
                        12'b011111010_001: ratio = -(24'b00000000_1111000011000000);
                        12'b011111010_100: ratio = -(24'b00000000_1111000101010000);
                        12'b011111010_111: ratio = -(24'b00000000_1111000111011110);
                        12'b011111011_010: ratio = -(24'b00000000_1111001001101010);
                        12'b011111011_101: ratio = -(24'b00000000_1111001011110010);
                        12'b011111100_000: ratio = -(24'b00000000_1111001101111000);
                        12'b011111100_011: ratio = -(24'b00000000_1111001111111011);
                        12'b011111100_110: ratio = -(24'b00000000_1111010001111100);
                        12'b011111101_001: ratio = -(24'b00000000_1111010011111010);
                        12'b011111101_100: ratio = -(24'b00000000_1111010101110101);
                        12'b011111101_111: ratio = -(24'b00000000_1111010111101101);
                        12'b011111110_010: ratio = -(24'b00000000_1111011001100011);
                        12'b011111110_101: ratio = -(24'b00000000_1111011011010110);
                        12'b011111111_000: ratio = -(24'b00000000_1111011101000110);
                        12'b011111111_011: ratio = -(24'b00000000_1111011110110100);
                        12'b011111111_110: ratio = -(24'b00000000_1111100000011111);
                        12'b100000000_001: ratio = -(24'b00000000_1111100010000111);
                        12'b100000000_100: ratio = -(24'b00000000_1111100011101101);
                        12'b100000000_111: ratio = -(24'b00000000_1111100101010000);
                        12'b100000001_010: ratio = -(24'b00000000_1111100110110000);
                        12'b100000001_101: ratio = -(24'b00000000_1111101000001101);
                        12'b100000010_000: ratio = -(24'b00000000_1111101001100111);
                        12'b100000010_011: ratio = -(24'b00000000_1111101010111111);
                        12'b100000010_110: ratio = -(24'b00000000_1111101100010100);
                        12'b100000011_001: ratio = -(24'b00000000_1111101101100111);
                        12'b100000011_100: ratio = -(24'b00000000_1111101110110110);
                        12'b100000011_111: ratio = -(24'b00000000_1111110000000011);
                        12'b100000100_010: ratio = -(24'b00000000_1111110001001101);
                        12'b100000100_101: ratio = -(24'b00000000_1111110010010100);
                        12'b100000101_000: ratio = -(24'b00000000_1111110011011001);
                        12'b100000101_011: ratio = -(24'b00000000_1111110100011010);
                        12'b100000101_110: ratio = -(24'b00000000_1111110101011001);
                        12'b100000110_001: ratio = -(24'b00000000_1111110110010101);
                        12'b100000110_100: ratio = -(24'b00000000_1111110111001111);
                        12'b100000110_111: ratio = -(24'b00000000_1111111000000101);
                        12'b100000111_010: ratio = -(24'b00000000_1111111000111001);
                        12'b100000111_101: ratio = -(24'b00000000_1111111001101010);
                        12'b100001000_000: ratio = -(24'b00000000_1111111010011000);
                        12'b100001000_011: ratio = -(24'b00000000_1111111011000100);
                        12'b100001000_110: ratio = -(24'b00000000_1111111011101101);
                        12'b100001001_001: ratio = -(24'b00000000_1111111100010010);
                        12'b100001001_100: ratio = -(24'b00000000_1111111100110101);
                        12'b100001001_111: ratio = -(24'b00000000_1111111101010110);
                        12'b100001010_010: ratio = -(24'b00000000_1111111101110011);
                        12'b100001010_101: ratio = -(24'b00000000_1111111110001110);
                        12'b100001011_000: ratio = -(24'b00000000_1111111110100110);
                        12'b100001011_011: ratio = -(24'b00000000_1111111110111011);
                        12'b100001011_110: ratio = -(24'b00000000_1111111111001101);
                        12'b100001100_001: ratio = -(24'b00000000_1111111111011100);
                        12'b100001100_100: ratio = -(24'b00000000_1111111111101001);
                        12'b100001100_111: ratio = -(24'b00000000_1111111111110011);
                        12'b100001101_010: ratio = -(24'b00000000_1111111111111010);
                        12'b100001101_101: ratio = -(24'b00000000_1111111111111110);
                        12'b100001110_000: ratio = -(24'b00000001_0000000000000000);
                        12'b100001110_011: ratio = -(24'b00000000_1111111111111110);
                        12'b100001110_110: ratio = -(24'b00000000_1111111111111010);
                        12'b100001111_001: ratio = -(24'b00000000_1111111111110011);
                        12'b100001111_100: ratio = -(24'b00000000_1111111111101001);
                        12'b100001111_111: ratio = -(24'b00000000_1111111111011100);
                        12'b100010000_010: ratio = -(24'b00000000_1111111111001101);
                        12'b100010000_101: ratio = -(24'b00000000_1111111110111011);
                        12'b100010001_000: ratio = -(24'b00000000_1111111110100110);
                        12'b100010001_011: ratio = -(24'b00000000_1111111110001110);
                        12'b100010001_110: ratio = -(24'b00000000_1111111101110011);
                        12'b100010010_001: ratio = -(24'b00000000_1111111101010110);
                        12'b100010010_100: ratio = -(24'b00000000_1111111100110101);
                        12'b100010010_111: ratio = -(24'b00000000_1111111100010010);
                        12'b100010011_010: ratio = -(24'b00000000_1111111011101101);
                        12'b100010011_101: ratio = -(24'b00000000_1111111011000100);
                        12'b100010100_000: ratio = -(24'b00000000_1111111010011000);
                        12'b100010100_011: ratio = -(24'b00000000_1111111001101010);
                        12'b100010100_110: ratio = -(24'b00000000_1111111000111001);
                        12'b100010101_001: ratio = -(24'b00000000_1111111000000101);
                        12'b100010101_100: ratio = -(24'b00000000_1111110111001111);
                        12'b100010101_111: ratio = -(24'b00000000_1111110110010101);
                        12'b100010110_010: ratio = -(24'b00000000_1111110101011001);
                        12'b100010110_101: ratio = -(24'b00000000_1111110100011010);
                        12'b100010111_000: ratio = -(24'b00000000_1111110011011001);
                        12'b100010111_011: ratio = -(24'b00000000_1111110010010100);
                        12'b100010111_110: ratio = -(24'b00000000_1111110001001101);
                        12'b100011000_001: ratio = -(24'b00000000_1111110000000011);
                        12'b100011000_100: ratio = -(24'b00000000_1111101110110110);
                        12'b100011000_111: ratio = -(24'b00000000_1111101101100111);
                        12'b100011001_010: ratio = -(24'b00000000_1111101100010100);
                        12'b100011001_101: ratio = -(24'b00000000_1111101010111111);
                        12'b100011010_000: ratio = -(24'b00000000_1111101001100111);
                        12'b100011010_011: ratio = -(24'b00000000_1111101000001101);
                        12'b100011010_110: ratio = -(24'b00000000_1111100110110000);
                        12'b100011011_001: ratio = -(24'b00000000_1111100101010000);
                        12'b100011011_100: ratio = -(24'b00000000_1111100011101101);
                        12'b100011011_111: ratio = -(24'b00000000_1111100010000111);
                        12'b100011100_010: ratio = -(24'b00000000_1111100000011111);
                        12'b100011100_101: ratio = -(24'b00000000_1111011110110100);
                        12'b100011101_000: ratio = -(24'b00000000_1111011101000110);
                        12'b100011101_011: ratio = -(24'b00000000_1111011011010110);
                        12'b100011101_110: ratio = -(24'b00000000_1111011001100011);
                        12'b100011110_001: ratio = -(24'b00000000_1111010111101101);
                        12'b100011110_100: ratio = -(24'b00000000_1111010101110101);
                        12'b100011110_111: ratio = -(24'b00000000_1111010011111010);
                        12'b100011111_010: ratio = -(24'b00000000_1111010001111100);
                        12'b100011111_101: ratio = -(24'b00000000_1111001111111011);
                        12'b100100000_000: ratio = -(24'b00000000_1111001101111000);
                        12'b100100000_011: ratio = -(24'b00000000_1111001011110010);
                        12'b100100000_110: ratio = -(24'b00000000_1111001001101010);
                        12'b100100001_001: ratio = -(24'b00000000_1111000111011110);
                        12'b100100001_100: ratio = -(24'b00000000_1111000101010000);
                        12'b100100001_111: ratio = -(24'b00000000_1111000011000000);
                        12'b100100010_010: ratio = -(24'b00000000_1111000000101101);
                        12'b100100010_101: ratio = -(24'b00000000_1110111110010111);
                        12'b100100011_000: ratio = -(24'b00000000_1110111011111111);
                        12'b100100011_011: ratio = -(24'b00000000_1110111001100100);
                        12'b100100011_110: ratio = -(24'b00000000_1110110111000110);
                        12'b100100100_001: ratio = -(24'b00000000_1110110100100110);
                        12'b100100100_100: ratio = -(24'b00000000_1110110010000011);
                        12'b100100100_111: ratio = -(24'b00000000_1110101111011101);
                        12'b100100101_010: ratio = -(24'b00000000_1110101100110101);
                        12'b100100101_101: ratio = -(24'b00000000_1110101010001011);
                        12'b100100110_000: ratio = -(24'b00000000_1110100111011110);
                        12'b100100110_011: ratio = -(24'b00000000_1110100100101110);
                        12'b100100110_110: ratio = -(24'b00000000_1110100001111100);
                        12'b100100111_001: ratio = -(24'b00000000_1110011111000111);
                        12'b100100111_100: ratio = -(24'b00000000_1110011100001111);
                        12'b100100111_111: ratio = -(24'b00000000_1110011001010101);
                        12'b100101000_010: ratio = -(24'b00000000_1110010110011001);
                        12'b100101000_101: ratio = -(24'b00000000_1110010011011010);
                        12'b100101001_000: ratio = -(24'b00000000_1110010000011001);
                        12'b100101001_011: ratio = -(24'b00000000_1110001101010101);
                        12'b100101001_110: ratio = -(24'b00000000_1110001010001110);
                        12'b100101010_001: ratio = -(24'b00000000_1110000111000101);
                        12'b100101010_100: ratio = -(24'b00000000_1110000011111010);
                        12'b100101010_111: ratio = -(24'b00000000_1110000000101100);
                        12'b100101011_010: ratio = -(24'b00000000_1101111101011011);
                        12'b100101011_101: ratio = -(24'b00000000_1101111010001001);
                        12'b100101100_000: ratio = -(24'b00000000_1101110110110011);
                        12'b100101100_011: ratio = -(24'b00000000_1101110011011100);
                        12'b100101100_110: ratio = -(24'b00000000_1101110000000010);
                        12'b100101101_001: ratio = -(24'b00000000_1101101100100101);
                        12'b100101101_100: ratio = -(24'b00000000_1101101001000110);
                        12'b100101101_111: ratio = -(24'b00000000_1101100101100101);
                        12'b100101110_010: ratio = -(24'b00000000_1101100010000001);
                        12'b100101110_101: ratio = -(24'b00000000_1101011110011011);
                        12'b100101111_000: ratio = -(24'b00000000_1101011010110011);
                        12'b100101111_011: ratio = -(24'b00000000_1101010111001000);
                        12'b100101111_110: ratio = -(24'b00000000_1101010011011011);
                        12'b100110000_001: ratio = -(24'b00000000_1101001111101011);
                        12'b100110000_100: ratio = -(24'b00000000_1101001011111001);
                        12'b100110000_111: ratio = -(24'b00000000_1101001000000101);
                        12'b100110001_010: ratio = -(24'b00000000_1101000100001111);
                        12'b100110001_101: ratio = -(24'b00000000_1101000000010110);
                        12'b100110010_000: ratio = -(24'b00000000_1100111100011011);
                        12'b100110010_011: ratio = -(24'b00000000_1100111000011110);
                        12'b100110010_110: ratio = -(24'b00000000_1100110100011110);
                        12'b100110011_001: ratio = -(24'b00000000_1100110000011101);
                        12'b100110011_100: ratio = -(24'b00000000_1100101100011001);
                        12'b100110011_111: ratio = -(24'b00000000_1100101000010010);
                        12'b100110100_010: ratio = -(24'b00000000_1100100100001010);
                        12'b100110100_101: ratio = -(24'b00000000_1100011111111111);
                        12'b100110101_000: ratio = -(24'b00000000_1100011011110011);
                        12'b100110101_011: ratio = -(24'b00000000_1100010111100100);
                        12'b100110101_110: ratio = -(24'b00000000_1100010011010010);
                        12'b100110110_001: ratio = -(24'b00000000_1100001110111111);
                        12'b100110110_100: ratio = -(24'b00000000_1100001010101001);
                        12'b100110110_111: ratio = -(24'b00000000_1100000110010010);
                        12'b100110111_010: ratio = -(24'b00000000_1100000001111000);
                        12'b100110111_101: ratio = -(24'b00000000_1011111101011100);
                        12'b100111000_000: ratio = -(24'b00000000_1011111000111110);
                        12'b100111000_011: ratio = -(24'b00000000_1011110100011110);
                        12'b100111000_110: ratio = -(24'b00000000_1011101111111100);
                        12'b100111001_001: ratio = -(24'b00000000_1011101011011000);
                        12'b100111001_100: ratio = -(24'b00000000_1011100110110010);
                        12'b100111001_111: ratio = -(24'b00000000_1011100010001001);
                        12'b100111010_010: ratio = -(24'b00000000_1011011101011111);
                        12'b100111010_101: ratio = -(24'b00000000_1011011000110011);
                        12'b100111011_000: ratio = -(24'b00000000_1011010100000100);
                        12'b100111011_011: ratio = -(24'b00000000_1011001111010100);
                        12'b100111011_110: ratio = -(24'b00000000_1011001010100010);
                        12'b100111100_001: ratio = -(24'b00000000_1011000101101110);
                        12'b100111100_100: ratio = -(24'b00000000_1011000000111000);
                        12'b100111100_111: ratio = -(24'b00000000_1010111011111111);
                        12'b100111101_010: ratio = -(24'b00000000_1010110111000101);
                        12'b100111101_101: ratio = -(24'b00000000_1010110010001001);
                        12'b100111110_000: ratio = -(24'b00000000_1010101101001100);
                        12'b100111110_011: ratio = -(24'b00000000_1010101000001100);
                        12'b100111110_110: ratio = -(24'b00000000_1010100011001010);
                        12'b100111111_001: ratio = -(24'b00000000_1010011110000111);
                        12'b100111111_100: ratio = -(24'b00000000_1010011001000010);
                        12'b100111111_111: ratio = -(24'b00000000_1010010011111011);
                        12'b101000000_010: ratio = -(24'b00000000_1010001110110010);
                        12'b101000000_101: ratio = -(24'b00000000_1010001001100111);
                        12'b101000001_000: ratio = -(24'b00000000_1010000100011011);
                        12'b101000001_011: ratio = -(24'b00000000_1001111111001100);
                        12'b101000001_110: ratio = -(24'b00000000_1001111001111100);
                        12'b101000010_001: ratio = -(24'b00000000_1001110100101011);
                        12'b101000010_100: ratio = -(24'b00000000_1001101111010111);
                        12'b101000010_111: ratio = -(24'b00000000_1001101010000010);
                        12'b101000011_010: ratio = -(24'b00000000_1001100100101011);
                        12'b101000011_101: ratio = -(24'b00000000_1001011111010011);
                        12'b101000100_000: ratio = -(24'b00000000_1001011001111001);
                        12'b101000100_011: ratio = -(24'b00000000_1001010100011101);
                        12'b101000100_110: ratio = -(24'b00000000_1001001110111111);
                        12'b101000101_001: ratio = -(24'b00000000_1001001001100000);
                        12'b101000101_100: ratio = -(24'b00000000_1001000011111111);
                        12'b101000101_111: ratio = -(24'b00000000_1000111110011101);
                        12'b101000110_010: ratio = -(24'b00000000_1000111000111001);
                        12'b101000110_101: ratio = -(24'b00000000_1000110011010100);
                        12'b101000111_000: ratio = -(24'b00000000_1000101101101101);
                        12'b101000111_011: ratio = -(24'b00000000_1000101000000100);
                        12'b101000111_110: ratio = -(24'b00000000_1000100010011010);
                        12'b101001000_001: ratio = -(24'b00000000_1000011100101111);
                        12'b101001000_100: ratio = -(24'b00000000_1000010111000010);
                        12'b101001000_111: ratio = -(24'b00000000_1000010001010100);
                        12'b101001001_010: ratio = -(24'b00000000_1000001011100100);
                        12'b101001001_101: ratio = -(24'b00000000_1000000101110010);
                        12'b101001010_000: ratio = -(24'b00000000_0111111111111111);
                        12'b101001010_011: ratio = -(24'b00000000_0111111010001011);
                        12'b101001010_110: ratio = -(24'b00000000_0111110100010110);
                        12'b101001011_001: ratio = -(24'b00000000_0111101110011111);
                        12'b101001011_100: ratio = -(24'b00000000_0111101000100111);
                        12'b101001011_111: ratio = -(24'b00000000_0111100010101101);
                        12'b101001100_010: ratio = -(24'b00000000_0111011100110010);
                        12'b101001100_101: ratio = -(24'b00000000_0111010110110110);
                        12'b101001101_000: ratio = -(24'b00000000_0111010000111000);
                        12'b101001101_011: ratio = -(24'b00000000_0111001010111001);
                        12'b101001101_110: ratio = -(24'b00000000_0111000100111001);
                        12'b101001110_001: ratio = -(24'b00000000_0110111110111000);
                        12'b101001110_100: ratio = -(24'b00000000_0110111000110101);
                        12'b101001110_111: ratio = -(24'b00000000_0110110010110010);
                        12'b101001111_010: ratio = -(24'b00000000_0110101100101101);
                        12'b101001111_101: ratio = -(24'b00000000_0110100110100111);
                        12'b101010000_000: ratio = -(24'b00000000_0110100000011111);
                        12'b101010000_011: ratio = -(24'b00000000_0110011010010111);
                        12'b101010000_110: ratio = -(24'b00000000_0110010100001101);
                        12'b101010001_001: ratio = -(24'b00000000_0110001110000011);
                        12'b101010001_100: ratio = -(24'b00000000_0110000111110111);
                        12'b101010001_111: ratio = -(24'b00000000_0110000001101010);
                        12'b101010010_010: ratio = -(24'b00000000_0101111011011100);
                        12'b101010010_101: ratio = -(24'b00000000_0101110101001101);
                        12'b101010011_000: ratio = -(24'b00000000_0101101110111110);
                        12'b101010011_011: ratio = -(24'b00000000_0101101000101101);
                        12'b101010011_110: ratio = -(24'b00000000_0101100010011011);
                        12'b101010100_001: ratio = -(24'b00000000_0101011100001000);
                        12'b101010100_100: ratio = -(24'b00000000_0101010101110100);
                        12'b101010100_111: ratio = -(24'b00000000_0101001111011111);
                        12'b101010101_010: ratio = -(24'b00000000_0101001001001001);
                        12'b101010101_101: ratio = -(24'b00000000_0101000010110011);
                        12'b101010110_000: ratio = -(24'b00000000_0100111100011011);
                        12'b101010110_011: ratio = -(24'b00000000_0100110110000011);
                        12'b101010110_110: ratio = -(24'b00000000_0100101111101010);
                        12'b101010111_001: ratio = -(24'b00000000_0100101001010000);
                        12'b101010111_100: ratio = -(24'b00000000_0100100010110101);
                        12'b101010111_111: ratio = -(24'b00000000_0100011100011001);
                        12'b101011000_010: ratio = -(24'b00000000_0100010101111101);
                        12'b101011000_101: ratio = -(24'b00000000_0100001111011111);
                        12'b101011001_000: ratio = -(24'b00000000_0100001001000001);
                        12'b101011001_011: ratio = -(24'b00000000_0100000010100011);
                        12'b101011001_110: ratio = -(24'b00000000_0011111100000011);
                        12'b101011010_001: ratio = -(24'b00000000_0011110101100011);
                        12'b101011010_100: ratio = -(24'b00000000_0011101111000011);
                        12'b101011010_111: ratio = -(24'b00000000_0011101000100001);
                        12'b101011011_010: ratio = -(24'b00000000_0011100001111111);
                        12'b101011011_101: ratio = -(24'b00000000_0011011011011100);
                        12'b101011100_000: ratio = -(24'b00000000_0011010100111001);
                        12'b101011100_011: ratio = -(24'b00000000_0011001110010101);
                        12'b101011100_110: ratio = -(24'b00000000_0011000111110001);
                        12'b101011101_001: ratio = -(24'b00000000_0011000001001100);
                        12'b101011101_100: ratio = -(24'b00000000_0010111010100110);
                        12'b101011101_111: ratio = -(24'b00000000_0010110100000000);
                        12'b101011110_010: ratio = -(24'b00000000_0010101101011010);
                        12'b101011110_101: ratio = -(24'b00000000_0010100110110011);
                        12'b101011111_000: ratio = -(24'b00000000_0010100000001100);
                        12'b101011111_011: ratio = -(24'b00000000_0010011001100100);
                        12'b101011111_110: ratio = -(24'b00000000_0010010010111011);
                        12'b101100000_001: ratio = -(24'b00000000_0010001100010011);
                        12'b101100000_100: ratio = -(24'b00000000_0010000101101010);
                        12'b101100000_111: ratio = -(24'b00000000_0001111111000000);
                        12'b101100001_010: ratio = -(24'b00000000_0001111000010110);
                        12'b101100001_101: ratio = -(24'b00000000_0001110001101100);
                        12'b101100010_000: ratio = -(24'b00000000_0001101011000010);
                        12'b101100010_011: ratio = -(24'b00000000_0001100100010111);
                        12'b101100010_110: ratio = -(24'b00000000_0001011101101100);
                        12'b101100011_001: ratio = -(24'b00000000_0001010111000001);
                        12'b101100011_100: ratio = -(24'b00000000_0001010000010101);
                        12'b101100011_111: ratio = -(24'b00000000_0001001001101010);
                        12'b101100100_010: ratio = -(24'b00000000_0001000010111110);
                        12'b101100100_101: ratio = -(24'b00000000_0000111100010010);
                        12'b101100101_000: ratio = -(24'b00000000_0000110101100101);
                        12'b101100101_011: ratio = -(24'b00000000_0000101110111001);
                        12'b101100101_110: ratio = -(24'b00000000_0000101000001100);
                        12'b101100110_001: ratio = -(24'b00000000_0000100001100000);
                        12'b101100110_100: ratio = -(24'b00000000_0000011010110011);
                        12'b101100110_111: ratio = -(24'b00000000_0000010100000110);
                        12'b101100111_010: ratio = -(24'b00000000_0000001101011001);
                        12'b101100111_101: ratio = -(24'b00000000_0000000110101100);
                        default: ratio = 24'b0;
                endcase
        end
endmodule

